module nivel
(
	input wire clk,rst,salto,
	input wire [9:0] hcount, vcount,
	input wire [9:0] origen_x,
	input wire [9:0] origen_y,
    output wire [3:0] rgb_out
);

// cambiar el tamaño segun la imagen
parameter tamano = 10'd64;
parameter y_tamano = 10'd64;
//parameter origen_x = 10'd200;
//reg[9:0] origen_x;
//parameter origen_y = 10'd200;

wire [12:0] lectura;
reg [3:0] w_rgb;
reg [2:0] registros [0:4095];



initial
begin
registros[0]= 3'b111;  
registros[1]= 3'b111;  
registros[2]= 3'b111;  
registros[3]= 3'b111;  
registros[4]= 3'b111;  
registros[5]= 3'b111;  
registros[6]= 3'b111;  
registros[7]= 3'b111;  
registros[8]= 3'b111;  
registros[9]= 3'b111;  
registros[10]= 3'b111;  
registros[11]= 3'b111;  
registros[12]= 3'b111;  
registros[13]= 3'b111;  
registros[14]= 3'b111;  
registros[15]= 3'b111;  
registros[16]= 3'b111;  
registros[17]= 3'b111;  
registros[18]= 3'b111;  
registros[19]= 3'b111;  
registros[20]= 3'b111;  
registros[21]= 3'b111;  
registros[22]= 3'b111;  
registros[23]= 3'b111;  
registros[24]= 3'b111;  
registros[25]= 3'b111;  
registros[26]= 3'b111;  
registros[27]= 3'b111;  
registros[28]= 3'b111;  
registros[29]= 3'b111;  
registros[30]= 3'b111;  
registros[31]= 3'b111;  
registros[32]= 3'b111;  
registros[33]= 3'b111;  
registros[34]= 3'b111;  
registros[35]= 3'b111;  
registros[36]= 3'b111;  
registros[37]= 3'b111;  
registros[38]= 3'b111;  
registros[39]= 3'b111;  
registros[40]= 3'b111;  
registros[41]= 3'b111;  
registros[42]= 3'b111;  
registros[43]= 3'b111;  
registros[44]= 3'b111;  
registros[45]= 3'b111;  
registros[46]= 3'b111;  
registros[47]= 3'b111;  
registros[48]= 3'b111;  
registros[49]= 3'b111;  
registros[50]= 3'b111;  
registros[51]= 3'b111;  
registros[52]= 3'b111;  
registros[53]= 3'b111;  
registros[54]= 3'b111;  
registros[55]= 3'b111;  
registros[56]= 3'b111;  
registros[57]= 3'b111;  
registros[58]= 3'b111;  
registros[59]= 3'b111;  
registros[60]= 3'b111;  
registros[61]= 3'b111;  
registros[62]= 3'b111;  
registros[63]= 3'b111;  
registros[64]= 3'b111;  
registros[65]= 3'b111;  
registros[66]= 3'b111;  
registros[67]= 3'b111;  
registros[68]= 3'b111;  
registros[69]= 3'b111;  
registros[70]= 3'b111;  
registros[71]= 3'b111;  
registros[72]= 3'b111;  
registros[73]= 3'b111;  
registros[74]= 3'b111;  
registros[75]= 3'b111;  
registros[76]= 3'b111;  
registros[77]= 3'b111;  
registros[78]= 3'b111;  
registros[79]= 3'b111;  
registros[80]= 3'b111;  
registros[81]= 3'b111;  
registros[82]= 3'b111;  
registros[83]= 3'b111;  
registros[84]= 3'b111;  
registros[85]= 3'b111;  
registros[86]= 3'b111;  
registros[87]= 3'b111;  
registros[88]= 3'b111;  
registros[89]= 3'b111;  
registros[90]= 3'b111;  
registros[91]= 3'b111;  
registros[92]= 3'b000;  
registros[93]= 3'b000;  
registros[94]= 3'b000;  
registros[95]= 3'b000;  
registros[96]= 3'b000;  
registros[97]= 3'b000;  
registros[98]= 3'b000;  
registros[99]= 3'b000;  
registros[100]= 3'b111;  
registros[101]= 3'b111;  
registros[102]= 3'b111;  
registros[103]= 3'b111;  
registros[104]= 3'b111;  
registros[105]= 3'b111;  
registros[106]= 3'b111;  
registros[107]= 3'b111;  
registros[108]= 3'b111;  
registros[109]= 3'b111;  
registros[110]= 3'b111;  
registros[111]= 3'b111;  
registros[112]= 3'b111;  
registros[113]= 3'b111;  
registros[114]= 3'b111;  
registros[115]= 3'b111;  
registros[116]= 3'b111;  
registros[117]= 3'b111;  
registros[118]= 3'b111;  
registros[119]= 3'b111;  
registros[120]= 3'b111;  
registros[121]= 3'b111;  
registros[122]= 3'b111;  
registros[123]= 3'b111;  
registros[124]= 3'b111;  
registros[125]= 3'b111;  
registros[126]= 3'b111;  
registros[127]= 3'b111;  
registros[128]= 3'b111;  
registros[129]= 3'b111;  
registros[130]= 3'b111;  
registros[131]= 3'b111;  
registros[132]= 3'b111;  
registros[133]= 3'b111;  
registros[134]= 3'b111;  
registros[135]= 3'b111;  
registros[136]= 3'b111;  
registros[137]= 3'b111;  
registros[138]= 3'b111;  
registros[139]= 3'b111;  
registros[140]= 3'b111;  
registros[141]= 3'b111;  
registros[142]= 3'b111;  
registros[143]= 3'b111;  
registros[144]= 3'b111;  
registros[145]= 3'b111;  
registros[146]= 3'b111;  
registros[147]= 3'b111;  
registros[148]= 3'b111;  
registros[149]= 3'b111;  
registros[150]= 3'b111;  
registros[151]= 3'b111;  
registros[152]= 3'b111;  
registros[153]= 3'b111;  
registros[154]= 3'b111;  
registros[155]= 3'b000;  
registros[156]= 3'b000;  
registros[157]= 3'b100;  
registros[158]= 3'b100;  
registros[159]= 3'b000;  
registros[160]= 3'b000;  
registros[161]= 3'b000;  
registros[162]= 3'b000;  
registros[163]= 3'b000;  
registros[164]= 3'b000;  
registros[165]= 3'b000;  
registros[166]= 3'b111;  
registros[167]= 3'b111;  
registros[168]= 3'b111;  
registros[169]= 3'b111;  
registros[170]= 3'b111;  
registros[171]= 3'b111;  
registros[172]= 3'b111;  
registros[173]= 3'b111;  
registros[174]= 3'b111;  
registros[175]= 3'b111;  
registros[176]= 3'b111;  
registros[177]= 3'b111;  
registros[178]= 3'b111;  
registros[179]= 3'b111;  
registros[180]= 3'b111;  
registros[181]= 3'b111;  
registros[182]= 3'b111;  
registros[183]= 3'b111;  
registros[184]= 3'b111;  
registros[185]= 3'b111;  
registros[186]= 3'b111;  
registros[187]= 3'b111;  
registros[188]= 3'b111;  
registros[189]= 3'b111;  
registros[190]= 3'b111;  
registros[191]= 3'b111;  
registros[192]= 3'b111;  
registros[193]= 3'b111;  
registros[194]= 3'b111;  
registros[195]= 3'b111;  
registros[196]= 3'b111;  
registros[197]= 3'b111;  
registros[198]= 3'b111;  
registros[199]= 3'b111;  
registros[200]= 3'b111;  
registros[201]= 3'b111;  
registros[202]= 3'b111;  
registros[203]= 3'b111;  
registros[204]= 3'b111;  
registros[205]= 3'b111;  
registros[206]= 3'b111;  
registros[207]= 3'b111;  
registros[208]= 3'b111;  
registros[209]= 3'b111;  
registros[210]= 3'b111;  
registros[211]= 3'b111;  
registros[212]= 3'b111;  
registros[213]= 3'b111;  
registros[214]= 3'b111;  
registros[215]= 3'b111;  
registros[216]= 3'b111;  
registros[217]= 3'b111;  
registros[218]= 3'b000;  
registros[219]= 3'b000;  
registros[220]= 3'b100;  
registros[221]= 3'b100;  
registros[222]= 3'b100;  
registros[223]= 3'b100;  
registros[224]= 3'b100;  
registros[225]= 3'b000;  
registros[226]= 3'b000;  
registros[227]= 3'b000;  
registros[228]= 3'b000;  
registros[229]= 3'b000;  
registros[230]= 3'b000;  
registros[231]= 3'b111;  
registros[232]= 3'b111;  
registros[233]= 3'b111;  
registros[234]= 3'b111;  
registros[235]= 3'b111;  
registros[236]= 3'b111;  
registros[237]= 3'b111;  
registros[238]= 3'b111;  
registros[239]= 3'b111;  
registros[240]= 3'b111;  
registros[241]= 3'b111;  
registros[242]= 3'b111;  
registros[243]= 3'b111;  
registros[244]= 3'b111;  
registros[245]= 3'b111;  
registros[246]= 3'b111;  
registros[247]= 3'b111;  
registros[248]= 3'b111;  
registros[249]= 3'b111;  
registros[250]= 3'b111;  
registros[251]= 3'b111;  
registros[252]= 3'b111;  
registros[253]= 3'b111;  
registros[254]= 3'b111;  
registros[255]= 3'b111;  
registros[256]= 3'b111;  
registros[257]= 3'b111;  
registros[258]= 3'b111;  
registros[259]= 3'b111;  
registros[260]= 3'b111;  
registros[261]= 3'b111;  
registros[262]= 3'b111;  
registros[263]= 3'b111;  
registros[264]= 3'b111;  
registros[265]= 3'b111;  
registros[266]= 3'b111;  
registros[267]= 3'b111;  
registros[268]= 3'b111;  
registros[269]= 3'b111;  
registros[270]= 3'b111;  
registros[271]= 3'b111;  
registros[272]= 3'b111;  
registros[273]= 3'b111;  
registros[274]= 3'b111;  
registros[275]= 3'b111;  
registros[276]= 3'b111;  
registros[277]= 3'b111;  
registros[278]= 3'b000;  
registros[279]= 3'b000;  
registros[280]= 3'b100;  
registros[281]= 3'b100;  
registros[282]= 3'b100;  
registros[283]= 3'b100;  
registros[284]= 3'b100;  
registros[285]= 3'b100;  
registros[286]= 3'b100;  
registros[287]= 3'b100;  
registros[288]= 3'b100;  
registros[289]= 3'b100;  
registros[290]= 3'b100;  
registros[291]= 3'b100;  
registros[292]= 3'b100;  
registros[293]= 3'b000;  
registros[294]= 3'b000;  
registros[295]= 3'b000;  
registros[296]= 3'b111;  
registros[297]= 3'b111;  
registros[298]= 3'b111;  
registros[299]= 3'b111;  
registros[300]= 3'b111;  
registros[301]= 3'b111;  
registros[302]= 3'b111;  
registros[303]= 3'b111;  
registros[304]= 3'b111;  
registros[305]= 3'b111;  
registros[306]= 3'b111;  
registros[307]= 3'b111;  
registros[308]= 3'b111;  
registros[309]= 3'b111;  
registros[310]= 3'b111;  
registros[311]= 3'b111;  
registros[312]= 3'b111;  
registros[313]= 3'b111;  
registros[314]= 3'b111;  
registros[315]= 3'b111;  
registros[316]= 3'b111;  
registros[317]= 3'b111;  
registros[318]= 3'b111;  
registros[319]= 3'b111;  
registros[320]= 3'b111;  
registros[321]= 3'b111;  
registros[322]= 3'b111;  
registros[323]= 3'b111;  
registros[324]= 3'b111;  
registros[325]= 3'b111;  
registros[326]= 3'b111;  
registros[327]= 3'b111;  
registros[328]= 3'b111;  
registros[329]= 3'b111;  
registros[330]= 3'b111;  
registros[331]= 3'b111;  
registros[332]= 3'b111;  
registros[333]= 3'b111;  
registros[334]= 3'b111;  
registros[335]= 3'b111;  
registros[336]= 3'b111;  
registros[337]= 3'b111;  
registros[338]= 3'b111;  
registros[339]= 3'b111;  
registros[340]= 3'b111;  
registros[341]= 3'b000;  
registros[342]= 3'b100;  
registros[343]= 3'b100;  
registros[344]= 3'b100;  
registros[345]= 3'b100;  
registros[346]= 3'b100;  
registros[347]= 3'b100;  
registros[348]= 3'b100;  
registros[349]= 3'b100;  
registros[350]= 3'b100;  
registros[351]= 3'b100;  
registros[352]= 3'b100;  
registros[353]= 3'b100;  
registros[354]= 3'b100;  
registros[355]= 3'b100;  
registros[356]= 3'b100;  
registros[357]= 3'b100;  
registros[358]= 3'b000;  
registros[359]= 3'b000;  
registros[360]= 3'b000;  
registros[361]= 3'b111;  
registros[362]= 3'b111;  
registros[363]= 3'b111;  
registros[364]= 3'b111;  
registros[365]= 3'b111;  
registros[366]= 3'b111;  
registros[367]= 3'b111;  
registros[368]= 3'b111;  
registros[369]= 3'b111;  
registros[370]= 3'b111;  
registros[371]= 3'b111;  
registros[372]= 3'b111;  
registros[373]= 3'b111;  
registros[374]= 3'b111;  
registros[375]= 3'b111;  
registros[376]= 3'b111;  
registros[377]= 3'b111;  
registros[378]= 3'b111;  
registros[379]= 3'b111;  
registros[380]= 3'b111;  
registros[381]= 3'b111;  
registros[382]= 3'b111;  
registros[383]= 3'b111;  
registros[384]= 3'b111;  
registros[385]= 3'b111;  
registros[386]= 3'b111;  
registros[387]= 3'b111;  
registros[388]= 3'b111;  
registros[389]= 3'b111;  
registros[390]= 3'b111;  
registros[391]= 3'b111;  
registros[392]= 3'b111;  
registros[393]= 3'b111;  
registros[394]= 3'b111;  
registros[395]= 3'b111;  
registros[396]= 3'b111;  
registros[397]= 3'b111;  
registros[398]= 3'b111;  
registros[399]= 3'b111;  
registros[400]= 3'b111;  
registros[401]= 3'b111;  
registros[402]= 3'b111;  
registros[403]= 3'b111;  
registros[404]= 3'b000;  
registros[405]= 3'b100;  
registros[406]= 3'b100;  
registros[407]= 3'b100;  
registros[408]= 3'b100;  
registros[409]= 3'b100;  
registros[410]= 3'b100;  
registros[411]= 3'b100;  
registros[412]= 3'b100;  
registros[413]= 3'b100;  
registros[414]= 3'b100;  
registros[415]= 3'b100;  
registros[416]= 3'b100;  
registros[417]= 3'b100;  
registros[418]= 3'b100;  
registros[419]= 3'b100;  
registros[420]= 3'b100;  
registros[421]= 3'b100;  
registros[422]= 3'b000;  
registros[423]= 3'b000;  
registros[424]= 3'b000;  
registros[425]= 3'b000;  
registros[426]= 3'b111;  
registros[427]= 3'b111;  
registros[428]= 3'b111;  
registros[429]= 3'b111;  
registros[430]= 3'b111;  
registros[431]= 3'b111;  
registros[432]= 3'b000;  
registros[433]= 3'b000;  
registros[434]= 3'b000;  
registros[435]= 3'b111;  
registros[436]= 3'b111;  
registros[437]= 3'b111;  
registros[438]= 3'b111;  
registros[439]= 3'b111;  
registros[440]= 3'b111;  
registros[441]= 3'b111;  
registros[442]= 3'b111;  
registros[443]= 3'b111;  
registros[444]= 3'b111;  
registros[445]= 3'b111;  
registros[446]= 3'b111;  
registros[447]= 3'b111;  
registros[448]= 3'b111;  
registros[449]= 3'b111;  
registros[450]= 3'b111;  
registros[451]= 3'b111;  
registros[452]= 3'b111;  
registros[453]= 3'b111;  
registros[454]= 3'b111;  
registros[455]= 3'b111;  
registros[456]= 3'b111;  
registros[457]= 3'b111;  
registros[458]= 3'b111;  
registros[459]= 3'b111;  
registros[460]= 3'b111;  
registros[461]= 3'b111;  
registros[462]= 3'b111;  
registros[463]= 3'b111;  
registros[464]= 3'b111;  
registros[465]= 3'b111;  
registros[466]= 3'b111;  
registros[467]= 3'b111;  
registros[468]= 3'b000;  
registros[469]= 3'b100;  
registros[470]= 3'b100;  
registros[471]= 3'b100;  
registros[472]= 3'b100;  
registros[473]= 3'b100;  
registros[474]= 3'b100;  
registros[475]= 3'b100;  
registros[476]= 3'b100;  
registros[477]= 3'b100;  
registros[478]= 3'b100;  
registros[479]= 3'b100;  
registros[480]= 3'b100;  
registros[481]= 3'b100;  
registros[482]= 3'b100;  
registros[483]= 3'b100;  
registros[484]= 3'b100;  
registros[485]= 3'b000;  
registros[486]= 3'b000;  
registros[487]= 3'b000;  
registros[488]= 3'b000;  
registros[489]= 3'b000;  
registros[490]= 3'b000;  
registros[491]= 3'b000;  
registros[492]= 3'b000;  
registros[493]= 3'b000;  
registros[494]= 3'b000;  
registros[495]= 3'b000;  
registros[496]= 3'b000;  
registros[497]= 3'b000;  
registros[498]= 3'b000;  
registros[499]= 3'b000;  
registros[500]= 3'b111;  
registros[501]= 3'b111;  
registros[502]= 3'b111;  
registros[503]= 3'b111;  
registros[504]= 3'b111;  
registros[505]= 3'b111;  
registros[506]= 3'b111;  
registros[507]= 3'b111;  
registros[508]= 3'b111;  
registros[509]= 3'b111;  
registros[510]= 3'b111;  
registros[511]= 3'b111;  
registros[512]= 3'b111;  
registros[513]= 3'b111;  
registros[514]= 3'b111;  
registros[515]= 3'b111;  
registros[516]= 3'b111;  
registros[517]= 3'b111;  
registros[518]= 3'b111;  
registros[519]= 3'b111;  
registros[520]= 3'b111;  
registros[521]= 3'b111;  
registros[522]= 3'b111;  
registros[523]= 3'b111;  
registros[524]= 3'b111;  
registros[525]= 3'b111;  
registros[526]= 3'b111;  
registros[527]= 3'b111;  
registros[528]= 3'b111;  
registros[529]= 3'b111;  
registros[530]= 3'b000;  
registros[531]= 3'b000;  
registros[532]= 3'b100;  
registros[533]= 3'b000;  
registros[534]= 3'b000;  
registros[535]= 3'b100;  
registros[536]= 3'b100;  
registros[537]= 3'b100;  
registros[538]= 3'b100;  
registros[539]= 3'b100;  
registros[540]= 3'b100;  
registros[541]= 3'b100;  
registros[542]= 3'b110;  
registros[543]= 3'b110;  
registros[544]= 3'b100;  
registros[545]= 3'b100;  
registros[546]= 3'b100;  
registros[547]= 3'b100;  
registros[548]= 3'b100;  
registros[549]= 3'b000;  
registros[550]= 3'b100;  
registros[551]= 3'b000;  
registros[552]= 3'b000;  
registros[553]= 3'b000;  
registros[554]= 3'b000;  
registros[555]= 3'b000;  
registros[556]= 3'b000;  
registros[557]= 3'b000;  
registros[558]= 3'b000;  
registros[559]= 3'b000;  
registros[560]= 3'b000;  
registros[561]= 3'b000;  
registros[562]= 3'b000;  
registros[563]= 3'b000;  
registros[564]= 3'b000;  
registros[565]= 3'b111;  
registros[566]= 3'b111;  
registros[567]= 3'b111;  
registros[568]= 3'b111;  
registros[569]= 3'b111;  
registros[570]= 3'b111;  
registros[571]= 3'b111;  
registros[572]= 3'b111;  
registros[573]= 3'b111;  
registros[574]= 3'b111;  
registros[575]= 3'b111;  
registros[576]= 3'b111;  
registros[577]= 3'b111;  
registros[578]= 3'b111;  
registros[579]= 3'b111;  
registros[580]= 3'b111;  
registros[581]= 3'b111;  
registros[582]= 3'b111;  
registros[583]= 3'b111;  
registros[584]= 3'b111;  
registros[585]= 3'b111;  
registros[586]= 3'b111;  
registros[587]= 3'b111;  
registros[588]= 3'b000;  
registros[589]= 3'b000;  
registros[590]= 3'b000;  
registros[591]= 3'b000;  
registros[592]= 3'b000;  
registros[593]= 3'b000;  
registros[594]= 3'b000;  
registros[595]= 3'b000;  
registros[596]= 3'b100;  
registros[597]= 3'b100;  
registros[598]= 3'b100;  
registros[599]= 3'b100;  
registros[600]= 3'b100;  
registros[601]= 3'b100;  
registros[602]= 3'b100;  
registros[603]= 3'b100;  
registros[604]= 3'b100;  
registros[605]= 3'b110;  
registros[606]= 3'b110;  
registros[607]= 3'b100;  
registros[608]= 3'b100;  
registros[609]= 3'b100;  
registros[610]= 3'b100;  
registros[611]= 3'b000;  
registros[612]= 3'b000;  
registros[613]= 3'b000;  
registros[614]= 3'b000;  
registros[615]= 3'b000;  
registros[616]= 3'b000;  
registros[617]= 3'b000;  
registros[618]= 3'b000;  
registros[619]= 3'b000;  
registros[620]= 3'b000;  
registros[621]= 3'b000;  
registros[622]= 3'b000;  
registros[623]= 3'b000;  
registros[624]= 3'b000;  
registros[625]= 3'b000;  
registros[626]= 3'b000;  
registros[627]= 3'b000;  
registros[628]= 3'b000;  
registros[629]= 3'b111;  
registros[630]= 3'b111;  
registros[631]= 3'b111;  
registros[632]= 3'b111;  
registros[633]= 3'b111;  
registros[634]= 3'b111;  
registros[635]= 3'b111;  
registros[636]= 3'b111;  
registros[637]= 3'b111;  
registros[638]= 3'b111;  
registros[639]= 3'b111;  
registros[640]= 3'b111;  
registros[641]= 3'b111;  
registros[642]= 3'b111;  
registros[643]= 3'b111;  
registros[644]= 3'b111;  
registros[645]= 3'b111;  
registros[646]= 3'b111;  
registros[647]= 3'b111;  
registros[648]= 3'b111;  
registros[649]= 3'b111;  
registros[650]= 3'b111;  
registros[651]= 3'b000;  
registros[652]= 3'b000;  
registros[653]= 3'b000;  
registros[654]= 3'b000;  
registros[655]= 3'b000;  
registros[656]= 3'b000;  
registros[657]= 3'b000;  
registros[658]= 3'b000;  
registros[659]= 3'b000;  
registros[660]= 3'b100;  
registros[661]= 3'b100;  
registros[662]= 3'b100;  
registros[663]= 3'b100;  
registros[664]= 3'b100;  
registros[665]= 3'b100;  
registros[666]= 3'b100;  
registros[667]= 3'b100;  
registros[668]= 3'b110;  
registros[669]= 3'b110;  
registros[670]= 3'b110;  
registros[671]= 3'b100;  
registros[672]= 3'b100;  
registros[673]= 3'b100;  
registros[674]= 3'b100;  
registros[675]= 3'b000;  
registros[676]= 3'b000;  
registros[677]= 3'b000;  
registros[678]= 3'b000;  
registros[679]= 3'b100;  
registros[680]= 3'b100;  
registros[681]= 3'b000;  
registros[682]= 3'b000;  
registros[683]= 3'b000;  
registros[684]= 3'b100;  
registros[685]= 3'b100;  
registros[686]= 3'b100;  
registros[687]= 3'b100;  
registros[688]= 3'b100;  
registros[689]= 3'b000;  
registros[690]= 3'b000;  
registros[691]= 3'b000;  
registros[692]= 3'b000;  
registros[693]= 3'b111;  
registros[694]= 3'b111;  
registros[695]= 3'b111;  
registros[696]= 3'b111;  
registros[697]= 3'b111;  
registros[698]= 3'b111;  
registros[699]= 3'b111;  
registros[700]= 3'b111;  
registros[701]= 3'b111;  
registros[702]= 3'b111;  
registros[703]= 3'b111;  
registros[704]= 3'b111;  
registros[705]= 3'b111;  
registros[706]= 3'b111;  
registros[707]= 3'b111;  
registros[708]= 3'b111;  
registros[709]= 3'b111;  
registros[710]= 3'b111;  
registros[711]= 3'b111;  
registros[712]= 3'b111;  
registros[713]= 3'b000;  
registros[714]= 3'b000;  
registros[715]= 3'b000;  
registros[716]= 3'b000;  
registros[717]= 3'b000;  
registros[718]= 3'b000;  
registros[719]= 3'b000;  
registros[720]= 3'b000;  
registros[721]= 3'b100;  
registros[722]= 3'b100;  
registros[723]= 3'b000;  
registros[724]= 3'b100;  
registros[725]= 3'b100;  
registros[726]= 3'b100;  
registros[727]= 3'b100;  
registros[728]= 3'b100;  
registros[729]= 3'b100;  
registros[730]= 3'b100;  
registros[731]= 3'b100;  
registros[732]= 3'b110;  
registros[733]= 3'b110;  
registros[734]= 3'b100;  
registros[735]= 3'b100;  
registros[736]= 3'b100;  
registros[737]= 3'b100;  
registros[738]= 3'b100;  
registros[739]= 3'b100;  
registros[740]= 3'b000;  
registros[741]= 3'b100;  
registros[742]= 3'b100;  
registros[743]= 3'b100;  
registros[744]= 3'b100;  
registros[745]= 3'b000;  
registros[746]= 3'b000;  
registros[747]= 3'b000;  
registros[748]= 3'b100;  
registros[749]= 3'b100;  
registros[750]= 3'b100;  
registros[751]= 3'b100;  
registros[752]= 3'b100;  
registros[753]= 3'b100;  
registros[754]= 3'b000;  
registros[755]= 3'b000;  
registros[756]= 3'b000;  
registros[757]= 3'b000;  
registros[758]= 3'b111;  
registros[759]= 3'b111;  
registros[760]= 3'b111;  
registros[761]= 3'b111;  
registros[762]= 3'b111;  
registros[763]= 3'b111;  
registros[764]= 3'b111;  
registros[765]= 3'b111;  
registros[766]= 3'b111;  
registros[767]= 3'b111;  
registros[768]= 3'b111;  
registros[769]= 3'b111;  
registros[770]= 3'b111;  
registros[771]= 3'b111;  
registros[772]= 3'b111;  
registros[773]= 3'b111;  
registros[774]= 3'b111;  
registros[775]= 3'b111;  
registros[776]= 3'b111;  
registros[777]= 3'b000;  
registros[778]= 3'b000;  
registros[779]= 3'b000;  
registros[780]= 3'b000;  
registros[781]= 3'b100;  
registros[782]= 3'b100;  
registros[783]= 3'b100;  
registros[784]= 3'b100;  
registros[785]= 3'b100;  
registros[786]= 3'b100;  
registros[787]= 3'b100;  
registros[788]= 3'b100;  
registros[789]= 3'b100;  
registros[790]= 3'b100;  
registros[791]= 3'b100;  
registros[792]= 3'b100;  
registros[793]= 3'b100;  
registros[794]= 3'b100;  
registros[795]= 3'b100;  
registros[796]= 3'b100;  
registros[797]= 3'b100;  
registros[798]= 3'b100;  
registros[799]= 3'b100;  
registros[800]= 3'b100;  
registros[801]= 3'b100;  
registros[802]= 3'b100;  
registros[803]= 3'b100;  
registros[804]= 3'b100;  
registros[805]= 3'b100;  
registros[806]= 3'b100;  
registros[807]= 3'b100;  
registros[808]= 3'b100;  
registros[809]= 3'b100;  
registros[810]= 3'b100;  
registros[811]= 3'b100;  
registros[812]= 3'b100;  
registros[813]= 3'b100;  
registros[814]= 3'b100;  
registros[815]= 3'b100;  
registros[816]= 3'b100;  
registros[817]= 3'b100;  
registros[818]= 3'b000;  
registros[819]= 3'b000;  
registros[820]= 3'b000;  
registros[821]= 3'b000;  
registros[822]= 3'b111;  
registros[823]= 3'b111;  
registros[824]= 3'b111;  
registros[825]= 3'b111;  
registros[826]= 3'b111;  
registros[827]= 3'b111;  
registros[828]= 3'b111;  
registros[829]= 3'b111;  
registros[830]= 3'b111;  
registros[831]= 3'b111;  
registros[832]= 3'b111;  
registros[833]= 3'b111;  
registros[834]= 3'b111;  
registros[835]= 3'b111;  
registros[836]= 3'b111;  
registros[837]= 3'b111;  
registros[838]= 3'b111;  
registros[839]= 3'b111;  
registros[840]= 3'b000;  
registros[841]= 3'b000;  
registros[842]= 3'b000;  
registros[843]= 3'b100;  
registros[844]= 3'b100;  
registros[845]= 3'b100;  
registros[846]= 3'b100;  
registros[847]= 3'b100;  
registros[848]= 3'b100;  
registros[849]= 3'b100;  
registros[850]= 3'b100;  
registros[851]= 3'b100;  
registros[852]= 3'b100;  
registros[853]= 3'b100;  
registros[854]= 3'b100;  
registros[855]= 3'b100;  
registros[856]= 3'b100;  
registros[857]= 3'b100;  
registros[858]= 3'b110;  
registros[859]= 3'b100;  
registros[860]= 3'b100;  
registros[861]= 3'b100;  
registros[862]= 3'b100;  
registros[863]= 3'b100;  
registros[864]= 3'b100;  
registros[865]= 3'b100;  
registros[866]= 3'b100;  
registros[867]= 3'b100;  
registros[868]= 3'b100;  
registros[869]= 3'b100;  
registros[870]= 3'b100;  
registros[871]= 3'b100;  
registros[872]= 3'b100;  
registros[873]= 3'b100;  
registros[874]= 3'b100;  
registros[875]= 3'b100;  
registros[876]= 3'b100;  
registros[877]= 3'b100;  
registros[878]= 3'b100;  
registros[879]= 3'b100;  
registros[880]= 3'b100;  
registros[881]= 3'b100;  
registros[882]= 3'b000;  
registros[883]= 3'b000;  
registros[884]= 3'b000;  
registros[885]= 3'b000;  
registros[886]= 3'b111;  
registros[887]= 3'b111;  
registros[888]= 3'b111;  
registros[889]= 3'b111;  
registros[890]= 3'b111;  
registros[891]= 3'b111;  
registros[892]= 3'b111;  
registros[893]= 3'b111;  
registros[894]= 3'b111;  
registros[895]= 3'b111;  
registros[896]= 3'b111;  
registros[897]= 3'b111;  
registros[898]= 3'b111;  
registros[899]= 3'b111;  
registros[900]= 3'b111;  
registros[901]= 3'b111;  
registros[902]= 3'b111;  
registros[903]= 3'b111;  
registros[904]= 3'b000;  
registros[905]= 3'b000;  
registros[906]= 3'b100;  
registros[907]= 3'b100;  
registros[908]= 3'b100;  
registros[909]= 3'b100;  
registros[910]= 3'b100;  
registros[911]= 3'b100;  
registros[912]= 3'b100;  
registros[913]= 3'b000;  
registros[914]= 3'b000;  
registros[915]= 3'b100;  
registros[916]= 3'b100;  
registros[917]= 3'b100;  
registros[918]= 3'b100;  
registros[919]= 3'b100;  
registros[920]= 3'b100;  
registros[921]= 3'b110;  
registros[922]= 3'b110;  
registros[923]= 3'b100;  
registros[924]= 3'b100;  
registros[925]= 3'b100;  
registros[926]= 3'b100;  
registros[927]= 3'b100;  
registros[928]= 3'b100;  
registros[929]= 3'b100;  
registros[930]= 3'b100;  
registros[931]= 3'b100;  
registros[932]= 3'b100;  
registros[933]= 3'b100;  
registros[934]= 3'b100;  
registros[935]= 3'b100;  
registros[936]= 3'b100;  
registros[937]= 3'b100;  
registros[938]= 3'b100;  
registros[939]= 3'b100;  
registros[940]= 3'b100;  
registros[941]= 3'b100;  
registros[942]= 3'b100;  
registros[943]= 3'b100;  
registros[944]= 3'b100;  
registros[945]= 3'b100;  
registros[946]= 3'b000;  
registros[947]= 3'b000;  
registros[948]= 3'b000;  
registros[949]= 3'b000;  
registros[950]= 3'b000;  
registros[951]= 3'b000;  
registros[952]= 3'b111;  
registros[953]= 3'b111;  
registros[954]= 3'b111;  
registros[955]= 3'b111;  
registros[956]= 3'b111;  
registros[957]= 3'b111;  
registros[958]= 3'b111;  
registros[959]= 3'b111;  
registros[960]= 3'b111;  
registros[961]= 3'b111;  
registros[962]= 3'b111;  
registros[963]= 3'b111;  
registros[964]= 3'b111;  
registros[965]= 3'b111;  
registros[966]= 3'b111;  
registros[967]= 3'b000;  
registros[968]= 3'b000;  
registros[969]= 3'b000;  
registros[970]= 3'b000;  
registros[971]= 3'b100;  
registros[972]= 3'b100;  
registros[973]= 3'b100;  
registros[974]= 3'b100;  
registros[975]= 3'b100;  
registros[976]= 3'b000;  
registros[977]= 3'b000;  
registros[978]= 3'b000;  
registros[979]= 3'b100;  
registros[980]= 3'b100;  
registros[981]= 3'b100;  
registros[982]= 3'b100;  
registros[983]= 3'b110;  
registros[984]= 3'b110;  
registros[985]= 3'b110;  
registros[986]= 3'b110;  
registros[987]= 3'b110;  
registros[988]= 3'b100;  
registros[989]= 3'b100;  
registros[990]= 3'b100;  
registros[991]= 3'b100;  
registros[992]= 3'b100;  
registros[993]= 3'b100;  
registros[994]= 3'b100;  
registros[995]= 3'b100;  
registros[996]= 3'b100;  
registros[997]= 3'b100;  
registros[998]= 3'b100;  
registros[999]= 3'b100;  
registros[1000]= 3'b100;  
registros[1001]= 3'b100;  
registros[1002]= 3'b100;  
registros[1003]= 3'b100;  
registros[1004]= 3'b100;  
registros[1005]= 3'b100;  
registros[1006]= 3'b100;  
registros[1007]= 3'b100;  
registros[1008]= 3'b100;  
registros[1009]= 3'b000;  
registros[1010]= 3'b000;  
registros[1011]= 3'b000;  
registros[1012]= 3'b000;  
registros[1013]= 3'b000;  
registros[1014]= 3'b000;  
registros[1015]= 3'b000;  
registros[1016]= 3'b000;  
registros[1017]= 3'b111;  
registros[1018]= 3'b111;  
registros[1019]= 3'b111;  
registros[1020]= 3'b111;  
registros[1021]= 3'b111;  
registros[1022]= 3'b111;  
registros[1023]= 3'b111;  
registros[1024]= 3'b111;  
registros[1025]= 3'b111;  
registros[1026]= 3'b111;  
registros[1027]= 3'b111;  
registros[1028]= 3'b111;  
registros[1029]= 3'b111;  
registros[1030]= 3'b000;  
registros[1031]= 3'b100;  
registros[1032]= 3'b000;  
registros[1033]= 3'b000;  
registros[1034]= 3'b000;  
registros[1035]= 3'b100;  
registros[1036]= 3'b100;  
registros[1037]= 3'b100;  
registros[1038]= 3'b100;  
registros[1039]= 3'b100;  
registros[1040]= 3'b100;  
registros[1041]= 3'b100;  
registros[1042]= 3'b100;  
registros[1043]= 3'b100;  
registros[1044]= 3'b100;  
registros[1045]= 3'b110;  
registros[1046]= 3'b110;  
registros[1047]= 3'b110;  
registros[1048]= 3'b110;  
registros[1049]= 3'b110;  
registros[1050]= 3'b110;  
registros[1051]= 3'b110;  
registros[1052]= 3'b110;  
registros[1053]= 3'b110;  
registros[1054]= 3'b100;  
registros[1055]= 3'b110;  
registros[1056]= 3'b100;  
registros[1057]= 3'b100;  
registros[1058]= 3'b100;  
registros[1059]= 3'b100;  
registros[1060]= 3'b100;  
registros[1061]= 3'b100;  
registros[1062]= 3'b100;  
registros[1063]= 3'b100;  
registros[1064]= 3'b100;  
registros[1065]= 3'b100;  
registros[1066]= 3'b100;  
registros[1067]= 3'b100;  
registros[1068]= 3'b100;  
registros[1069]= 3'b100;  
registros[1070]= 3'b100;  
registros[1071]= 3'b000;  
registros[1072]= 3'b000;  
registros[1073]= 3'b000;  
registros[1074]= 3'b000;  
registros[1075]= 3'b000;  
registros[1076]= 3'b000;  
registros[1077]= 3'b000;  
registros[1078]= 3'b000;  
registros[1079]= 3'b000;  
registros[1080]= 3'b000;  
registros[1081]= 3'b111;  
registros[1082]= 3'b111;  
registros[1083]= 3'b111;  
registros[1084]= 3'b111;  
registros[1085]= 3'b111;  
registros[1086]= 3'b111;  
registros[1087]= 3'b111;  
registros[1088]= 3'b111;  
registros[1089]= 3'b111;  
registros[1090]= 3'b111;  
registros[1091]= 3'b111;  
registros[1092]= 3'b111;  
registros[1093]= 3'b000;  
registros[1094]= 3'b100;  
registros[1095]= 3'b100;  
registros[1096]= 3'b100;  
registros[1097]= 3'b100;  
registros[1098]= 3'b100;  
registros[1099]= 3'b100;  
registros[1100]= 3'b100;  
registros[1101]= 3'b100;  
registros[1102]= 3'b100;  
registros[1103]= 3'b100;  
registros[1104]= 3'b100;  
registros[1105]= 3'b100;  
registros[1106]= 3'b100;  
registros[1107]= 3'b100;  
registros[1108]= 3'b110;  
registros[1109]= 3'b110;  
registros[1110]= 3'b110;  
registros[1111]= 3'b110;  
registros[1112]= 3'b110;  
registros[1113]= 3'b110;  
registros[1114]= 3'b110;  
registros[1115]= 3'b110;  
registros[1116]= 3'b110;  
registros[1117]= 3'b100;  
registros[1118]= 3'b100;  
registros[1119]= 3'b100;  
registros[1120]= 3'b100;  
registros[1121]= 3'b100;  
registros[1122]= 3'b100;  
registros[1123]= 3'b100;  
registros[1124]= 3'b100;  
registros[1125]= 3'b100;  
registros[1126]= 3'b100;  
registros[1127]= 3'b100;  
registros[1128]= 3'b100;  
registros[1129]= 3'b100;  
registros[1130]= 3'b100;  
registros[1131]= 3'b100;  
registros[1132]= 3'b100;  
registros[1133]= 3'b000;  
registros[1134]= 3'b000;  
registros[1135]= 3'b000;  
registros[1136]= 3'b000;  
registros[1137]= 3'b000;  
registros[1138]= 3'b000;  
registros[1139]= 3'b000;  
registros[1140]= 3'b000;  
registros[1141]= 3'b000;  
registros[1142]= 3'b000;  
registros[1143]= 3'b000;  
registros[1144]= 3'b000;  
registros[1145]= 3'b000;  
registros[1146]= 3'b111;  
registros[1147]= 3'b111;  
registros[1148]= 3'b111;  
registros[1149]= 3'b111;  
registros[1150]= 3'b111;  
registros[1151]= 3'b111;  
registros[1152]= 3'b111;  
registros[1153]= 3'b111;  
registros[1154]= 3'b111;  
registros[1155]= 3'b111;  
registros[1156]= 3'b000;  
registros[1157]= 3'b100;  
registros[1158]= 3'b000;  
registros[1159]= 3'b100;  
registros[1160]= 3'b100;  
registros[1161]= 3'b100;  
registros[1162]= 3'b100;  
registros[1163]= 3'b100;  
registros[1164]= 3'b100;  
registros[1165]= 3'b100;  
registros[1166]= 3'b100;  
registros[1167]= 3'b100;  
registros[1168]= 3'b100;  
registros[1169]= 3'b110;  
registros[1170]= 3'b100;  
registros[1171]= 3'b100;  
registros[1172]= 3'b110;  
registros[1173]= 3'b110;  
registros[1174]= 3'b110;  
registros[1175]= 3'b110;  
registros[1176]= 3'b110;  
registros[1177]= 3'b110;  
registros[1178]= 3'b110;  
registros[1179]= 3'b110;  
registros[1180]= 3'b100;  
registros[1181]= 3'b100;  
registros[1182]= 3'b100;  
registros[1183]= 3'b110;  
registros[1184]= 3'b100;  
registros[1185]= 3'b100;  
registros[1186]= 3'b100;  
registros[1187]= 3'b100;  
registros[1188]= 3'b100;  
registros[1189]= 3'b100;  
registros[1190]= 3'b100;  
registros[1191]= 3'b100;  
registros[1192]= 3'b100;  
registros[1193]= 3'b100;  
registros[1194]= 3'b100;  
registros[1195]= 3'b100;  
registros[1196]= 3'b000;  
registros[1197]= 3'b000;  
registros[1198]= 3'b000;  
registros[1199]= 3'b000;  
registros[1200]= 3'b000;  
registros[1201]= 3'b000;  
registros[1202]= 3'b000;  
registros[1203]= 3'b000;  
registros[1204]= 3'b000;  
registros[1205]= 3'b000;  
registros[1206]= 3'b000;  
registros[1207]= 3'b000;  
registros[1208]= 3'b000;  
registros[1209]= 3'b000;  
registros[1210]= 3'b000;  
registros[1211]= 3'b111;  
registros[1212]= 3'b111;  
registros[1213]= 3'b111;  
registros[1214]= 3'b111;  
registros[1215]= 3'b111;  
registros[1216]= 3'b111;  
registros[1217]= 3'b111;  
registros[1218]= 3'b111;  
registros[1219]= 3'b000;  
registros[1220]= 3'b000;  
registros[1221]= 3'b000;  
registros[1222]= 3'b100;  
registros[1223]= 3'b100;  
registros[1224]= 3'b100;  
registros[1225]= 3'b100;  
registros[1226]= 3'b100;  
registros[1227]= 3'b100;  
registros[1228]= 3'b100;  
registros[1229]= 3'b100;  
registros[1230]= 3'b100;  
registros[1231]= 3'b100;  
registros[1232]= 3'b100;  
registros[1233]= 3'b100;  
registros[1234]= 3'b110;  
registros[1235]= 3'b100;  
registros[1236]= 3'b100;  
registros[1237]= 3'b110;  
registros[1238]= 3'b110;  
registros[1239]= 3'b110;  
registros[1240]= 3'b110;  
registros[1241]= 3'b110;  
registros[1242]= 3'b110;  
registros[1243]= 3'b100;  
registros[1244]= 3'b100;  
registros[1245]= 3'b100;  
registros[1246]= 3'b100;  
registros[1247]= 3'b100;  
registros[1248]= 3'b100;  
registros[1249]= 3'b100;  
registros[1250]= 3'b100;  
registros[1251]= 3'b100;  
registros[1252]= 3'b100;  
registros[1253]= 3'b100;  
registros[1254]= 3'b100;  
registros[1255]= 3'b100;  
registros[1256]= 3'b100;  
registros[1257]= 3'b100;  
registros[1258]= 3'b000;  
registros[1259]= 3'b000;  
registros[1260]= 3'b000;  
registros[1261]= 3'b000;  
registros[1262]= 3'b000;  
registros[1263]= 3'b000;  
registros[1264]= 3'b000;  
registros[1265]= 3'b000;  
registros[1266]= 3'b000;  
registros[1267]= 3'b000;  
registros[1268]= 3'b000;  
registros[1269]= 3'b000;  
registros[1270]= 3'b000;  
registros[1271]= 3'b000;  
registros[1272]= 3'b000;  
registros[1273]= 3'b000;  
registros[1274]= 3'b000;  
registros[1275]= 3'b111;  
registros[1276]= 3'b111;  
registros[1277]= 3'b111;  
registros[1278]= 3'b111;  
registros[1279]= 3'b111;  
registros[1280]= 3'b111;  
registros[1281]= 3'b111;  
registros[1282]= 3'b111;  
registros[1283]= 3'b000;  
registros[1284]= 3'b000;  
registros[1285]= 3'b100;  
registros[1286]= 3'b100;  
registros[1287]= 3'b100;  
registros[1288]= 3'b100;  
registros[1289]= 3'b100;  
registros[1290]= 3'b100;  
registros[1291]= 3'b100;  
registros[1292]= 3'b100;  
registros[1293]= 3'b100;  
registros[1294]= 3'b100;  
registros[1295]= 3'b100;  
registros[1296]= 3'b100;  
registros[1297]= 3'b100;  
registros[1298]= 3'b100;  
registros[1299]= 3'b100;  
registros[1300]= 3'b100;  
registros[1301]= 3'b110;  
registros[1302]= 3'b110;  
registros[1303]= 3'b110;  
registros[1304]= 3'b110;  
registros[1305]= 3'b110;  
registros[1306]= 3'b100;  
registros[1307]= 3'b110;  
registros[1308]= 3'b110;  
registros[1309]= 3'b110;  
registros[1310]= 3'b100;  
registros[1311]= 3'b100;  
registros[1312]= 3'b100;  
registros[1313]= 3'b100;  
registros[1314]= 3'b100;  
registros[1315]= 3'b100;  
registros[1316]= 3'b100;  
registros[1317]= 3'b100;  
registros[1318]= 3'b100;  
registros[1319]= 3'b100;  
registros[1320]= 3'b100;  
registros[1321]= 3'b000;  
registros[1322]= 3'b000;  
registros[1323]= 3'b000;  
registros[1324]= 3'b000;  
registros[1325]= 3'b000;  
registros[1326]= 3'b000;  
registros[1327]= 3'b000;  
registros[1328]= 3'b000;  
registros[1329]= 3'b000;  
registros[1330]= 3'b000;  
registros[1331]= 3'b000;  
registros[1332]= 3'b000;  
registros[1333]= 3'b000;  
registros[1334]= 3'b000;  
registros[1335]= 3'b000;  
registros[1336]= 3'b000;  
registros[1337]= 3'b000;  
registros[1338]= 3'b000;  
registros[1339]= 3'b000;  
registros[1340]= 3'b111;  
registros[1341]= 3'b111;  
registros[1342]= 3'b111;  
registros[1343]= 3'b111;  
registros[1344]= 3'b111;  
registros[1345]= 3'b111;  
registros[1346]= 3'b000;  
registros[1347]= 3'b100;  
registros[1348]= 3'b100;  
registros[1349]= 3'b100;  
registros[1350]= 3'b100;  
registros[1351]= 3'b100;  
registros[1352]= 3'b100;  
registros[1353]= 3'b100;  
registros[1354]= 3'b100;  
registros[1355]= 3'b100;  
registros[1356]= 3'b100;  
registros[1357]= 3'b100;  
registros[1358]= 3'b100;  
registros[1359]= 3'b100;  
registros[1360]= 3'b100;  
registros[1361]= 3'b100;  
registros[1362]= 3'b100;  
registros[1363]= 3'b100;  
registros[1364]= 3'b100;  
registros[1365]= 3'b100;  
registros[1366]= 3'b110;  
registros[1367]= 3'b110;  
registros[1368]= 3'b100;  
registros[1369]= 3'b100;  
registros[1370]= 3'b110;  
registros[1371]= 3'b110;  
registros[1372]= 3'b110;  
registros[1373]= 3'b110;  
registros[1374]= 3'b110;  
registros[1375]= 3'b100;  
registros[1376]= 3'b100;  
registros[1377]= 3'b100;  
registros[1378]= 3'b100;  
registros[1379]= 3'b100;  
registros[1380]= 3'b100;  
registros[1381]= 3'b100;  
registros[1382]= 3'b100;  
registros[1383]= 3'b100;  
registros[1384]= 3'b100;  
registros[1385]= 3'b000;  
registros[1386]= 3'b000;  
registros[1387]= 3'b000;  
registros[1388]= 3'b000;  
registros[1389]= 3'b000;  
registros[1390]= 3'b000;  
registros[1391]= 3'b000;  
registros[1392]= 3'b000;  
registros[1393]= 3'b000;  
registros[1394]= 3'b000;  
registros[1395]= 3'b000;  
registros[1396]= 3'b000;  
registros[1397]= 3'b000;  
registros[1398]= 3'b000;  
registros[1399]= 3'b000;  
registros[1400]= 3'b000;  
registros[1401]= 3'b000;  
registros[1402]= 3'b000;  
registros[1403]= 3'b000;  
registros[1404]= 3'b000;  
registros[1405]= 3'b111;  
registros[1406]= 3'b111;  
registros[1407]= 3'b111;  
registros[1408]= 3'b111;  
registros[1409]= 3'b000;  
registros[1410]= 3'b100;  
registros[1411]= 3'b100;  
registros[1412]= 3'b100;  
registros[1413]= 3'b100;  
registros[1414]= 3'b100;  
registros[1415]= 3'b100;  
registros[1416]= 3'b100;  
registros[1417]= 3'b100;  
registros[1418]= 3'b100;  
registros[1419]= 3'b100;  
registros[1420]= 3'b100;  
registros[1421]= 3'b100;  
registros[1422]= 3'b100;  
registros[1423]= 3'b100;  
registros[1424]= 3'b100;  
registros[1425]= 3'b100;  
registros[1426]= 3'b100;  
registros[1427]= 3'b100;  
registros[1428]= 3'b100;  
registros[1429]= 3'b100;  
registros[1430]= 3'b100;  
registros[1431]= 3'b100;  
registros[1432]= 3'b100;  
registros[1433]= 3'b110;  
registros[1434]= 3'b110;  
registros[1435]= 3'b110;  
registros[1436]= 3'b110;  
registros[1437]= 3'b110;  
registros[1438]= 3'b110;  
registros[1439]= 3'b110;  
registros[1440]= 3'b100;  
registros[1441]= 3'b100;  
registros[1442]= 3'b100;  
registros[1443]= 3'b100;  
registros[1444]= 3'b100;  
registros[1445]= 3'b100;  
registros[1446]= 3'b100;  
registros[1447]= 3'b100;  
registros[1448]= 3'b100;  
registros[1449]= 3'b100;  
registros[1450]= 3'b000;  
registros[1451]= 3'b000;  
registros[1452]= 3'b000;  
registros[1453]= 3'b000;  
registros[1454]= 3'b000;  
registros[1455]= 3'b000;  
registros[1456]= 3'b000;  
registros[1457]= 3'b000;  
registros[1458]= 3'b000;  
registros[1459]= 3'b000;  
registros[1460]= 3'b000;  
registros[1461]= 3'b000;  
registros[1462]= 3'b000;  
registros[1463]= 3'b000;  
registros[1464]= 3'b000;  
registros[1465]= 3'b000;  
registros[1466]= 3'b000;  
registros[1467]= 3'b000;  
registros[1468]= 3'b000;  
registros[1469]= 3'b000;  
registros[1470]= 3'b111;  
registros[1471]= 3'b111;  
registros[1472]= 3'b111;  
registros[1473]= 3'b100;  
registros[1474]= 3'b100;  
registros[1475]= 3'b100;  
registros[1476]= 3'b100;  
registros[1477]= 3'b100;  
registros[1478]= 3'b100;  
registros[1479]= 3'b100;  
registros[1480]= 3'b100;  
registros[1481]= 3'b100;  
registros[1482]= 3'b100;  
registros[1483]= 3'b100;  
registros[1484]= 3'b100;  
registros[1485]= 3'b100;  
registros[1486]= 3'b100;  
registros[1487]= 3'b100;  
registros[1488]= 3'b100;  
registros[1489]= 3'b100;  
registros[1490]= 3'b100;  
registros[1491]= 3'b110;  
registros[1492]= 3'b110;  
registros[1493]= 3'b110;  
registros[1494]= 3'b100;  
registros[1495]= 3'b100;  
registros[1496]= 3'b100;  
registros[1497]= 3'b110;  
registros[1498]= 3'b110;  
registros[1499]= 3'b110;  
registros[1500]= 3'b110;  
registros[1501]= 3'b110;  
registros[1502]= 3'b110;  
registros[1503]= 3'b110;  
registros[1504]= 3'b100;  
registros[1505]= 3'b100;  
registros[1506]= 3'b100;  
registros[1507]= 3'b100;  
registros[1508]= 3'b100;  
registros[1509]= 3'b100;  
registros[1510]= 3'b100;  
registros[1511]= 3'b100;  
registros[1512]= 3'b100;  
registros[1513]= 3'b100;  
registros[1514]= 3'b100;  
registros[1515]= 3'b100;  
registros[1516]= 3'b100;  
registros[1517]= 3'b000;  
registros[1518]= 3'b000;  
registros[1519]= 3'b000;  
registros[1520]= 3'b000;  
registros[1521]= 3'b000;  
registros[1522]= 3'b000;  
registros[1523]= 3'b000;  
registros[1524]= 3'b000;  
registros[1525]= 3'b000;  
registros[1526]= 3'b000;  
registros[1527]= 3'b000;  
registros[1528]= 3'b000;  
registros[1529]= 3'b000;  
registros[1530]= 3'b000;  
registros[1531]= 3'b000;  
registros[1532]= 3'b000;  
registros[1533]= 3'b000;  
registros[1534]= 3'b111;  
registros[1535]= 3'b111;  
registros[1536]= 3'b000;  
registros[1537]= 3'b100;  
registros[1538]= 3'b100;  
registros[1539]= 3'b100;  
registros[1540]= 3'b100;  
registros[1541]= 3'b100;  
registros[1542]= 3'b100;  
registros[1543]= 3'b110;  
registros[1544]= 3'b110;  
registros[1545]= 3'b110;  
registros[1546]= 3'b110;  
registros[1547]= 3'b100;  
registros[1548]= 3'b100;  
registros[1549]= 3'b100;  
registros[1550]= 3'b100;  
registros[1551]= 3'b100;  
registros[1552]= 3'b100;  
registros[1553]= 3'b100;  
registros[1554]= 3'b100;  
registros[1555]= 3'b110;  
registros[1556]= 3'b110;  
registros[1557]= 3'b110;  
registros[1558]= 3'b100;  
registros[1559]= 3'b100;  
registros[1560]= 3'b100;  
registros[1561]= 3'b110;  
registros[1562]= 3'b110;  
registros[1563]= 3'b110;  
registros[1564]= 3'b110;  
registros[1565]= 3'b110;  
registros[1566]= 3'b110;  
registros[1567]= 3'b100;  
registros[1568]= 3'b100;  
registros[1569]= 3'b100;  
registros[1570]= 3'b100;  
registros[1571]= 3'b100;  
registros[1572]= 3'b100;  
registros[1573]= 3'b100;  
registros[1574]= 3'b100;  
registros[1575]= 3'b100;  
registros[1576]= 3'b100;  
registros[1577]= 3'b100;  
registros[1578]= 3'b100;  
registros[1579]= 3'b100;  
registros[1580]= 3'b100;  
registros[1581]= 3'b100;  
registros[1582]= 3'b000;  
registros[1583]= 3'b000;  
registros[1584]= 3'b000;  
registros[1585]= 3'b000;  
registros[1586]= 3'b000;  
registros[1587]= 3'b000;  
registros[1588]= 3'b000;  
registros[1589]= 3'b000;  
registros[1590]= 3'b000;  
registros[1591]= 3'b000;  
registros[1592]= 3'b000;  
registros[1593]= 3'b000;  
registros[1594]= 3'b000;  
registros[1595]= 3'b000;  
registros[1596]= 3'b000;  
registros[1597]= 3'b111;  
registros[1598]= 3'b111;  
registros[1599]= 3'b111;  
registros[1600]= 3'b000;  
registros[1601]= 3'b100;  
registros[1602]= 3'b100;  
registros[1603]= 3'b100;  
registros[1604]= 3'b100;  
registros[1605]= 3'b100;  
registros[1606]= 3'b100;  
registros[1607]= 3'b100;  
registros[1608]= 3'b110;  
registros[1609]= 3'b110;  
registros[1610]= 3'b110;  
registros[1611]= 3'b100;  
registros[1612]= 3'b100;  
registros[1613]= 3'b100;  
registros[1614]= 3'b100;  
registros[1615]= 3'b100;  
registros[1616]= 3'b100;  
registros[1617]= 3'b100;  
registros[1618]= 3'b110;  
registros[1619]= 3'b110;  
registros[1620]= 3'b110;  
registros[1621]= 3'b110;  
registros[1622]= 3'b110;  
registros[1623]= 3'b110;  
registros[1624]= 3'b100;  
registros[1625]= 3'b100;  
registros[1626]= 3'b110;  
registros[1627]= 3'b110;  
registros[1628]= 3'b110;  
registros[1629]= 3'b110;  
registros[1630]= 3'b100;  
registros[1631]= 3'b100;  
registros[1632]= 3'b100;  
registros[1633]= 3'b100;  
registros[1634]= 3'b100;  
registros[1635]= 3'b100;  
registros[1636]= 3'b100;  
registros[1637]= 3'b100;  
registros[1638]= 3'b100;  
registros[1639]= 3'b100;  
registros[1640]= 3'b100;  
registros[1641]= 3'b100;  
registros[1642]= 3'b100;  
registros[1643]= 3'b100;  
registros[1644]= 3'b100;  
registros[1645]= 3'b100;  
registros[1646]= 3'b100;  
registros[1647]= 3'b100;  
registros[1648]= 3'b100;  
registros[1649]= 3'b000;  
registros[1650]= 3'b000;  
registros[1651]= 3'b100;  
registros[1652]= 3'b000;  
registros[1653]= 3'b000;  
registros[1654]= 3'b000;  
registros[1655]= 3'b000;  
registros[1656]= 3'b000;  
registros[1657]= 3'b000;  
registros[1658]= 3'b000;  
registros[1659]= 3'b000;  
registros[1660]= 3'b111;  
registros[1661]= 3'b111;  
registros[1662]= 3'b111;  
registros[1663]= 3'b111;  
registros[1664]= 3'b111;  
registros[1665]= 3'b100;  
registros[1666]= 3'b100;  
registros[1667]= 3'b100;  
registros[1668]= 3'b100;  
registros[1669]= 3'b100;  
registros[1670]= 3'b100;  
registros[1671]= 3'b100;  
registros[1672]= 3'b110;  
registros[1673]= 3'b110;  
registros[1674]= 3'b100;  
registros[1675]= 3'b100;  
registros[1676]= 3'b100;  
registros[1677]= 3'b110;  
registros[1678]= 3'b110;  
registros[1679]= 3'b110;  
registros[1680]= 3'b110;  
registros[1681]= 3'b110;  
registros[1682]= 3'b110;  
registros[1683]= 3'b110;  
registros[1684]= 3'b110;  
registros[1685]= 3'b110;  
registros[1686]= 3'b110;  
registros[1687]= 3'b110;  
registros[1688]= 3'b100;  
registros[1689]= 3'b100;  
registros[1690]= 3'b100;  
registros[1691]= 3'b100;  
registros[1692]= 3'b100;  
registros[1693]= 3'b100;  
registros[1694]= 3'b100;  
registros[1695]= 3'b100;  
registros[1696]= 3'b100;  
registros[1697]= 3'b100;  
registros[1698]= 3'b100;  
registros[1699]= 3'b100;  
registros[1700]= 3'b100;  
registros[1701]= 3'b100;  
registros[1702]= 3'b100;  
registros[1703]= 3'b100;  
registros[1704]= 3'b100;  
registros[1705]= 3'b100;  
registros[1706]= 3'b100;  
registros[1707]= 3'b100;  
registros[1708]= 3'b100;  
registros[1709]= 3'b100;  
registros[1710]= 3'b100;  
registros[1711]= 3'b100;  
registros[1712]= 3'b100;  
registros[1713]= 3'b100;  
registros[1714]= 3'b100;  
registros[1715]= 3'b100;  
registros[1716]= 3'b100;  
registros[1717]= 3'b000;  
registros[1718]= 3'b000;  
registros[1719]= 3'b000;  
registros[1720]= 3'b000;  
registros[1721]= 3'b000;  
registros[1722]= 3'b000;  
registros[1723]= 3'b000;  
registros[1724]= 3'b111;  
registros[1725]= 3'b111;  
registros[1726]= 3'b111;  
registros[1727]= 3'b111;  
registros[1728]= 3'b111;  
registros[1729]= 3'b000;  
registros[1730]= 3'b100;  
registros[1731]= 3'b100;  
registros[1732]= 3'b100;  
registros[1733]= 3'b100;  
registros[1734]= 3'b100;  
registros[1735]= 3'b100;  
registros[1736]= 3'b100;  
registros[1737]= 3'b100;  
registros[1738]= 3'b100;  
registros[1739]= 3'b100;  
registros[1740]= 3'b100;  
registros[1741]= 3'b110;  
registros[1742]= 3'b110;  
registros[1743]= 3'b110;  
registros[1744]= 3'b110;  
registros[1745]= 3'b110;  
registros[1746]= 3'b110;  
registros[1747]= 3'b110;  
registros[1748]= 3'b110;  
registros[1749]= 3'b110;  
registros[1750]= 3'b110;  
registros[1751]= 3'b110;  
registros[1752]= 3'b110;  
registros[1753]= 3'b100;  
registros[1754]= 3'b100;  
registros[1755]= 3'b100;  
registros[1756]= 3'b100;  
registros[1757]= 3'b100;  
registros[1758]= 3'b100;  
registros[1759]= 3'b100;  
registros[1760]= 3'b100;  
registros[1761]= 3'b100;  
registros[1762]= 3'b100;  
registros[1763]= 3'b100;  
registros[1764]= 3'b100;  
registros[1765]= 3'b100;  
registros[1766]= 3'b100;  
registros[1767]= 3'b100;  
registros[1768]= 3'b100;  
registros[1769]= 3'b100;  
registros[1770]= 3'b100;  
registros[1771]= 3'b100;  
registros[1772]= 3'b100;  
registros[1773]= 3'b100;  
registros[1774]= 3'b000;  
registros[1775]= 3'b100;  
registros[1776]= 3'b100;  
registros[1777]= 3'b100;  
registros[1778]= 3'b100;  
registros[1779]= 3'b100;  
registros[1780]= 3'b100;  
registros[1781]= 3'b100;  
registros[1782]= 3'b100;  
registros[1783]= 3'b000;  
registros[1784]= 3'b000;  
registros[1785]= 3'b000;  
registros[1786]= 3'b000;  
registros[1787]= 3'b000;  
registros[1788]= 3'b000;  
registros[1789]= 3'b000;  
registros[1790]= 3'b111;  
registros[1791]= 3'b111;  
registros[1792]= 3'b111;  
registros[1793]= 3'b111;  
registros[1794]= 3'b100;  
registros[1795]= 3'b100;  
registros[1796]= 3'b100;  
registros[1797]= 3'b100;  
registros[1798]= 3'b100;  
registros[1799]= 3'b100;  
registros[1800]= 3'b100;  
registros[1801]= 3'b100;  
registros[1802]= 3'b110;  
registros[1803]= 3'b100;  
registros[1804]= 3'b100;  
registros[1805]= 3'b110;  
registros[1806]= 3'b110;  
registros[1807]= 3'b110;  
registros[1808]= 3'b110;  
registros[1809]= 3'b110;  
registros[1810]= 3'b110;  
registros[1811]= 3'b110;  
registros[1812]= 3'b110;  
registros[1813]= 3'b110;  
registros[1814]= 3'b110;  
registros[1815]= 3'b110;  
registros[1816]= 3'b110;  
registros[1817]= 3'b110;  
registros[1818]= 3'b100;  
registros[1819]= 3'b100;  
registros[1820]= 3'b100;  
registros[1821]= 3'b100;  
registros[1822]= 3'b100;  
registros[1823]= 3'b100;  
registros[1824]= 3'b100;  
registros[1825]= 3'b100;  
registros[1826]= 3'b100;  
registros[1827]= 3'b100;  
registros[1828]= 3'b110;  
registros[1829]= 3'b110;  
registros[1830]= 3'b100;  
registros[1831]= 3'b100;  
registros[1832]= 3'b100;  
registros[1833]= 3'b100;  
registros[1834]= 3'b100;  
registros[1835]= 3'b000;  
registros[1836]= 3'b000;  
registros[1837]= 3'b100;  
registros[1838]= 3'b100;  
registros[1839]= 3'b100;  
registros[1840]= 3'b100;  
registros[1841]= 3'b100;  
registros[1842]= 3'b100;  
registros[1843]= 3'b100;  
registros[1844]= 3'b100;  
registros[1845]= 3'b100;  
registros[1846]= 3'b100;  
registros[1847]= 3'b000;  
registros[1848]= 3'b000;  
registros[1849]= 3'b000;  
registros[1850]= 3'b000;  
registros[1851]= 3'b000;  
registros[1852]= 3'b000;  
registros[1853]= 3'b000;  
registros[1854]= 3'b000;  
registros[1855]= 3'b111;  
registros[1856]= 3'b111;  
registros[1857]= 3'b111;  
registros[1858]= 3'b100;  
registros[1859]= 3'b100;  
registros[1860]= 3'b100;  
registros[1861]= 3'b100;  
registros[1862]= 3'b100;  
registros[1863]= 3'b100;  
registros[1864]= 3'b100;  
registros[1865]= 3'b100;  
registros[1866]= 3'b110;  
registros[1867]= 3'b100;  
registros[1868]= 3'b110;  
registros[1869]= 3'b110;  
registros[1870]= 3'b110;  
registros[1871]= 3'b110;  
registros[1872]= 3'b110;  
registros[1873]= 3'b110;  
registros[1874]= 3'b110;  
registros[1875]= 3'b110;  
registros[1876]= 3'b110;  
registros[1877]= 3'b110;  
registros[1878]= 3'b110;  
registros[1879]= 3'b110;  
registros[1880]= 3'b110;  
registros[1881]= 3'b110;  
registros[1882]= 3'b100;  
registros[1883]= 3'b110;  
registros[1884]= 3'b110;  
registros[1885]= 3'b100;  
registros[1886]= 3'b100;  
registros[1887]= 3'b100;  
registros[1888]= 3'b100;  
registros[1889]= 3'b100;  
registros[1890]= 3'b100;  
registros[1891]= 3'b100;  
registros[1892]= 3'b100;  
registros[1893]= 3'b100;  
registros[1894]= 3'b110;  
registros[1895]= 3'b100;  
registros[1896]= 3'b100;  
registros[1897]= 3'b100;  
registros[1898]= 3'b100;  
registros[1899]= 3'b000;  
registros[1900]= 3'b100;  
registros[1901]= 3'b100;  
registros[1902]= 3'b100;  
registros[1903]= 3'b100;  
registros[1904]= 3'b100;  
registros[1905]= 3'b100;  
registros[1906]= 3'b100;  
registros[1907]= 3'b100;  
registros[1908]= 3'b100;  
registros[1909]= 3'b100;  
registros[1910]= 3'b000;  
registros[1911]= 3'b000;  
registros[1912]= 3'b000;  
registros[1913]= 3'b000;  
registros[1914]= 3'b000;  
registros[1915]= 3'b000;  
registros[1916]= 3'b000;  
registros[1917]= 3'b000;  
registros[1918]= 3'b000;  
registros[1919]= 3'b111;  
registros[1920]= 3'b111;  
registros[1921]= 3'b111;  
registros[1922]= 3'b100;  
registros[1923]= 3'b100;  
registros[1924]= 3'b100;  
registros[1925]= 3'b100;  
registros[1926]= 3'b100;  
registros[1927]= 3'b100;  
registros[1928]= 3'b100;  
registros[1929]= 3'b100;  
registros[1930]= 3'b100;  
registros[1931]= 3'b100;  
registros[1932]= 3'b110;  
registros[1933]= 3'b110;  
registros[1934]= 3'b110;  
registros[1935]= 3'b110;  
registros[1936]= 3'b110;  
registros[1937]= 3'b110;  
registros[1938]= 3'b110;  
registros[1939]= 3'b110;  
registros[1940]= 3'b110;  
registros[1941]= 3'b110;  
registros[1942]= 3'b110;  
registros[1943]= 3'b110;  
registros[1944]= 3'b110;  
registros[1945]= 3'b110;  
registros[1946]= 3'b110;  
registros[1947]= 3'b110;  
registros[1948]= 3'b110;  
registros[1949]= 3'b100;  
registros[1950]= 3'b100;  
registros[1951]= 3'b100;  
registros[1952]= 3'b110;  
registros[1953]= 3'b100;  
registros[1954]= 3'b100;  
registros[1955]= 3'b100;  
registros[1956]= 3'b100;  
registros[1957]= 3'b100;  
registros[1958]= 3'b100;  
registros[1959]= 3'b100;  
registros[1960]= 3'b100;  
registros[1961]= 3'b100;  
registros[1962]= 3'b100;  
registros[1963]= 3'b100;  
registros[1964]= 3'b100;  
registros[1965]= 3'b100;  
registros[1966]= 3'b100;  
registros[1967]= 3'b100;  
registros[1968]= 3'b100;  
registros[1969]= 3'b100;  
registros[1970]= 3'b100;  
registros[1971]= 3'b100;  
registros[1972]= 3'b100;  
registros[1973]= 3'b100;  
registros[1974]= 3'b000;  
registros[1975]= 3'b000;  
registros[1976]= 3'b000;  
registros[1977]= 3'b000;  
registros[1978]= 3'b000;  
registros[1979]= 3'b000;  
registros[1980]= 3'b000;  
registros[1981]= 3'b000;  
registros[1982]= 3'b000;  
registros[1983]= 3'b111;  
registros[1984]= 3'b111;  
registros[1985]= 3'b111;  
registros[1986]= 3'b100;  
registros[1987]= 3'b100;  
registros[1988]= 3'b100;  
registros[1989]= 3'b100;  
registros[1990]= 3'b100;  
registros[1991]= 3'b100;  
registros[1992]= 3'b100;  
registros[1993]= 3'b100;  
registros[1994]= 3'b100;  
registros[1995]= 3'b100;  
registros[1996]= 3'b110;  
registros[1997]= 3'b110;  
registros[1998]= 3'b110;  
registros[1999]= 3'b110;  
registros[2000]= 3'b110;  
registros[2001]= 3'b110;  
registros[2002]= 3'b110;  
registros[2003]= 3'b110;  
registros[2004]= 3'b110;  
registros[2005]= 3'b110;  
registros[2006]= 3'b110;  
registros[2007]= 3'b110;  
registros[2008]= 3'b110;  
registros[2009]= 3'b110;  
registros[2010]= 3'b110;  
registros[2011]= 3'b100;  
registros[2012]= 3'b100;  
registros[2013]= 3'b110;  
registros[2014]= 3'b100;  
registros[2015]= 3'b100;  
registros[2016]= 3'b110;  
registros[2017]= 3'b110;  
registros[2018]= 3'b110;  
registros[2019]= 3'b110;  
registros[2020]= 3'b100;  
registros[2021]= 3'b100;  
registros[2022]= 3'b100;  
registros[2023]= 3'b100;  
registros[2024]= 3'b100;  
registros[2025]= 3'b100;  
registros[2026]= 3'b100;  
registros[2027]= 3'b100;  
registros[2028]= 3'b100;  
registros[2029]= 3'b100;  
registros[2030]= 3'b100;  
registros[2031]= 3'b100;  
registros[2032]= 3'b100;  
registros[2033]= 3'b100;  
registros[2034]= 3'b100;  
registros[2035]= 3'b100;  
registros[2036]= 3'b100;  
registros[2037]= 3'b100;  
registros[2038]= 3'b000;  
registros[2039]= 3'b000;  
registros[2040]= 3'b000;  
registros[2041]= 3'b000;  
registros[2042]= 3'b000;  
registros[2043]= 3'b000;  
registros[2044]= 3'b000;  
registros[2045]= 3'b000;  
registros[2046]= 3'b000;  
registros[2047]= 3'b111;  
registros[2048]= 3'b111;  
registros[2049]= 3'b111;  
registros[2050]= 3'b100;  
registros[2051]= 3'b100;  
registros[2052]= 3'b100;  
registros[2053]= 3'b100;  
registros[2054]= 3'b100;  
registros[2055]= 3'b100;  
registros[2056]= 3'b100;  
registros[2057]= 3'b100;  
registros[2058]= 3'b100;  
registros[2059]= 3'b110;  
registros[2060]= 3'b110;  
registros[2061]= 3'b110;  
registros[2062]= 3'b110;  
registros[2063]= 3'b110;  
registros[2064]= 3'b110;  
registros[2065]= 3'b110;  
registros[2066]= 3'b110;  
registros[2067]= 3'b110;  
registros[2068]= 3'b110;  
registros[2069]= 3'b110;  
registros[2070]= 3'b110;  
registros[2071]= 3'b100;  
registros[2072]= 3'b100;  
registros[2073]= 3'b110;  
registros[2074]= 3'b110;  
registros[2075]= 3'b100;  
registros[2076]= 3'b100;  
registros[2077]= 3'b110;  
registros[2078]= 3'b110;  
registros[2079]= 3'b100;  
registros[2080]= 3'b100;  
registros[2081]= 3'b110;  
registros[2082]= 3'b110;  
registros[2083]= 3'b110;  
registros[2084]= 3'b100;  
registros[2085]= 3'b100;  
registros[2086]= 3'b100;  
registros[2087]= 3'b100;  
registros[2088]= 3'b100;  
registros[2089]= 3'b100;  
registros[2090]= 3'b100;  
registros[2091]= 3'b100;  
registros[2092]= 3'b100;  
registros[2093]= 3'b100;  
registros[2094]= 3'b100;  
registros[2095]= 3'b100;  
registros[2096]= 3'b100;  
registros[2097]= 3'b100;  
registros[2098]= 3'b100;  
registros[2099]= 3'b100;  
registros[2100]= 3'b100;  
registros[2101]= 3'b100;  
registros[2102]= 3'b000;  
registros[2103]= 3'b000;  
registros[2104]= 3'b000;  
registros[2105]= 3'b000;  
registros[2106]= 3'b000;  
registros[2107]= 3'b000;  
registros[2108]= 3'b000;  
registros[2109]= 3'b000;  
registros[2110]= 3'b000;  
registros[2111]= 3'b111;  
registros[2112]= 3'b111;  
registros[2113]= 3'b000;  
registros[2114]= 3'b100;  
registros[2115]= 3'b100;  
registros[2116]= 3'b100;  
registros[2117]= 3'b100;  
registros[2118]= 3'b110;  
registros[2119]= 3'b110;  
registros[2120]= 3'b110;  
registros[2121]= 3'b100;  
registros[2122]= 3'b100;  
registros[2123]= 3'b100;  
registros[2124]= 3'b110;  
registros[2125]= 3'b110;  
registros[2126]= 3'b110;  
registros[2127]= 3'b110;  
registros[2128]= 3'b110;  
registros[2129]= 3'b110;  
registros[2130]= 3'b110;  
registros[2131]= 3'b110;  
registros[2132]= 3'b110;  
registros[2133]= 3'b110;  
registros[2134]= 3'b100;  
registros[2135]= 3'b100;  
registros[2136]= 3'b100;  
registros[2137]= 3'b110;  
registros[2138]= 3'b110;  
registros[2139]= 3'b100;  
registros[2140]= 3'b100;  
registros[2141]= 3'b100;  
registros[2142]= 3'b100;  
registros[2143]= 3'b100;  
registros[2144]= 3'b100;  
registros[2145]= 3'b100;  
registros[2146]= 3'b100;  
registros[2147]= 3'b100;  
registros[2148]= 3'b100;  
registros[2149]= 3'b100;  
registros[2150]= 3'b100;  
registros[2151]= 3'b100;  
registros[2152]= 3'b100;  
registros[2153]= 3'b100;  
registros[2154]= 3'b100;  
registros[2155]= 3'b100;  
registros[2156]= 3'b100;  
registros[2157]= 3'b100;  
registros[2158]= 3'b100;  
registros[2159]= 3'b100;  
registros[2160]= 3'b100;  
registros[2161]= 3'b100;  
registros[2162]= 3'b100;  
registros[2163]= 3'b100;  
registros[2164]= 3'b100;  
registros[2165]= 3'b100;  
registros[2166]= 3'b100;  
registros[2167]= 3'b000;  
registros[2168]= 3'b000;  
registros[2169]= 3'b000;  
registros[2170]= 3'b000;  
registros[2171]= 3'b000;  
registros[2172]= 3'b000;  
registros[2173]= 3'b000;  
registros[2174]= 3'b000;  
registros[2175]= 3'b111;  
registros[2176]= 3'b111;  
registros[2177]= 3'b000;  
registros[2178]= 3'b100;  
registros[2179]= 3'b100;  
registros[2180]= 3'b110;  
registros[2181]= 3'b110;  
registros[2182]= 3'b110;  
registros[2183]= 3'b110;  
registros[2184]= 3'b110;  
registros[2185]= 3'b110;  
registros[2186]= 3'b100;  
registros[2187]= 3'b100;  
registros[2188]= 3'b100;  
registros[2189]= 3'b110;  
registros[2190]= 3'b110;  
registros[2191]= 3'b110;  
registros[2192]= 3'b110;  
registros[2193]= 3'b110;  
registros[2194]= 3'b110;  
registros[2195]= 3'b110;  
registros[2196]= 3'b100;  
registros[2197]= 3'b100;  
registros[2198]= 3'b100;  
registros[2199]= 3'b100;  
registros[2200]= 3'b100;  
registros[2201]= 3'b110;  
registros[2202]= 3'b110;  
registros[2203]= 3'b110;  
registros[2204]= 3'b110;  
registros[2205]= 3'b100;  
registros[2206]= 3'b100;  
registros[2207]= 3'b100;  
registros[2208]= 3'b100;  
registros[2209]= 3'b100;  
registros[2210]= 3'b100;  
registros[2211]= 3'b100;  
registros[2212]= 3'b100;  
registros[2213]= 3'b100;  
registros[2214]= 3'b100;  
registros[2215]= 3'b100;  
registros[2216]= 3'b100;  
registros[2217]= 3'b100;  
registros[2218]= 3'b100;  
registros[2219]= 3'b100;  
registros[2220]= 3'b100;  
registros[2221]= 3'b100;  
registros[2222]= 3'b100;  
registros[2223]= 3'b100;  
registros[2224]= 3'b100;  
registros[2225]= 3'b100;  
registros[2226]= 3'b100;  
registros[2227]= 3'b100;  
registros[2228]= 3'b100;  
registros[2229]= 3'b000;  
registros[2230]= 3'b000;  
registros[2231]= 3'b000;  
registros[2232]= 3'b000;  
registros[2233]= 3'b000;  
registros[2234]= 3'b000;  
registros[2235]= 3'b000;  
registros[2236]= 3'b000;  
registros[2237]= 3'b000;  
registros[2238]= 3'b000;  
registros[2239]= 3'b111;  
registros[2240]= 3'b111;  
registros[2241]= 3'b100;  
registros[2242]= 3'b100;  
registros[2243]= 3'b100;  
registros[2244]= 3'b110;  
registros[2245]= 3'b110;  
registros[2246]= 3'b110;  
registros[2247]= 3'b110;  
registros[2248]= 3'b110;  
registros[2249]= 3'b110;  
registros[2250]= 3'b110;  
registros[2251]= 3'b110;  
registros[2252]= 3'b100;  
registros[2253]= 3'b100;  
registros[2254]= 3'b110;  
registros[2255]= 3'b110;  
registros[2256]= 3'b110;  
registros[2257]= 3'b110;  
registros[2258]= 3'b100;  
registros[2259]= 3'b100;  
registros[2260]= 3'b100;  
registros[2261]= 3'b100;  
registros[2262]= 3'b100;  
registros[2263]= 3'b100;  
registros[2264]= 3'b100;  
registros[2265]= 3'b100;  
registros[2266]= 3'b110;  
registros[2267]= 3'b110;  
registros[2268]= 3'b110;  
registros[2269]= 3'b100;  
registros[2270]= 3'b100;  
registros[2271]= 3'b100;  
registros[2272]= 3'b100;  
registros[2273]= 3'b100;  
registros[2274]= 3'b100;  
registros[2275]= 3'b100;  
registros[2276]= 3'b100;  
registros[2277]= 3'b100;  
registros[2278]= 3'b100;  
registros[2279]= 3'b100;  
registros[2280]= 3'b100;  
registros[2281]= 3'b100;  
registros[2282]= 3'b100;  
registros[2283]= 3'b100;  
registros[2284]= 3'b100;  
registros[2285]= 3'b100;  
registros[2286]= 3'b100;  
registros[2287]= 3'b100;  
registros[2288]= 3'b100;  
registros[2289]= 3'b100;  
registros[2290]= 3'b100;  
registros[2291]= 3'b100;  
registros[2292]= 3'b100;  
registros[2293]= 3'b000;  
registros[2294]= 3'b000;  
registros[2295]= 3'b000;  
registros[2296]= 3'b000;  
registros[2297]= 3'b000;  
registros[2298]= 3'b000;  
registros[2299]= 3'b000;  
registros[2300]= 3'b000;  
registros[2301]= 3'b000;  
registros[2302]= 3'b000;  
registros[2303]= 3'b111;  
registros[2304]= 3'b000;  
registros[2305]= 3'b100;  
registros[2306]= 3'b100;  
registros[2307]= 3'b100;  
registros[2308]= 3'b100;  
registros[2309]= 3'b110;  
registros[2310]= 3'b110;  
registros[2311]= 3'b110;  
registros[2312]= 3'b110;  
registros[2313]= 3'b110;  
registros[2314]= 3'b110;  
registros[2315]= 3'b110;  
registros[2316]= 3'b110;  
registros[2317]= 3'b100;  
registros[2318]= 3'b100;  
registros[2319]= 3'b100;  
registros[2320]= 3'b100;  
registros[2321]= 3'b100;  
registros[2322]= 3'b100;  
registros[2323]= 3'b100;  
registros[2324]= 3'b100;  
registros[2325]= 3'b100;  
registros[2326]= 3'b100;  
registros[2327]= 3'b100;  
registros[2328]= 3'b100;  
registros[2329]= 3'b100;  
registros[2330]= 3'b100;  
registros[2331]= 3'b110;  
registros[2332]= 3'b110;  
registros[2333]= 3'b100;  
registros[2334]= 3'b100;  
registros[2335]= 3'b100;  
registros[2336]= 3'b100;  
registros[2337]= 3'b100;  
registros[2338]= 3'b100;  
registros[2339]= 3'b100;  
registros[2340]= 3'b100;  
registros[2341]= 3'b100;  
registros[2342]= 3'b100;  
registros[2343]= 3'b100;  
registros[2344]= 3'b100;  
registros[2345]= 3'b100;  
registros[2346]= 3'b100;  
registros[2347]= 3'b100;  
registros[2348]= 3'b100;  
registros[2349]= 3'b100;  
registros[2350]= 3'b100;  
registros[2351]= 3'b100;  
registros[2352]= 3'b100;  
registros[2353]= 3'b100;  
registros[2354]= 3'b100;  
registros[2355]= 3'b100;  
registros[2356]= 3'b100;  
registros[2357]= 3'b000;  
registros[2358]= 3'b000;  
registros[2359]= 3'b000;  
registros[2360]= 3'b000;  
registros[2361]= 3'b000;  
registros[2362]= 3'b000;  
registros[2363]= 3'b000;  
registros[2364]= 3'b000;  
registros[2365]= 3'b000;  
registros[2366]= 3'b000;  
registros[2367]= 3'b111;  
registros[2368]= 3'b000;  
registros[2369]= 3'b100;  
registros[2370]= 3'b100;  
registros[2371]= 3'b100;  
registros[2372]= 3'b100;  
registros[2373]= 3'b100;  
registros[2374]= 3'b110;  
registros[2375]= 3'b110;  
registros[2376]= 3'b110;  
registros[2377]= 3'b110;  
registros[2378]= 3'b100;  
registros[2379]= 3'b100;  
registros[2380]= 3'b100;  
registros[2381]= 3'b100;  
registros[2382]= 3'b100;  
registros[2383]= 3'b100;  
registros[2384]= 3'b100;  
registros[2385]= 3'b100;  
registros[2386]= 3'b100;  
registros[2387]= 3'b100;  
registros[2388]= 3'b100;  
registros[2389]= 3'b100;  
registros[2390]= 3'b100;  
registros[2391]= 3'b100;  
registros[2392]= 3'b100;  
registros[2393]= 3'b100;  
registros[2394]= 3'b100;  
registros[2395]= 3'b100;  
registros[2396]= 3'b100;  
registros[2397]= 3'b100;  
registros[2398]= 3'b100;  
registros[2399]= 3'b100;  
registros[2400]= 3'b100;  
registros[2401]= 3'b100;  
registros[2402]= 3'b100;  
registros[2403]= 3'b100;  
registros[2404]= 3'b100;  
registros[2405]= 3'b100;  
registros[2406]= 3'b100;  
registros[2407]= 3'b100;  
registros[2408]= 3'b100;  
registros[2409]= 3'b100;  
registros[2410]= 3'b100;  
registros[2411]= 3'b100;  
registros[2412]= 3'b100;  
registros[2413]= 3'b100;  
registros[2414]= 3'b100;  
registros[2415]= 3'b100;  
registros[2416]= 3'b100;  
registros[2417]= 3'b100;  
registros[2418]= 3'b100;  
registros[2419]= 3'b000;  
registros[2420]= 3'b000;  
registros[2421]= 3'b000;  
registros[2422]= 3'b000;  
registros[2423]= 3'b000;  
registros[2424]= 3'b000;  
registros[2425]= 3'b000;  
registros[2426]= 3'b000;  
registros[2427]= 3'b000;  
registros[2428]= 3'b000;  
registros[2429]= 3'b000;  
registros[2430]= 3'b000;  
registros[2431]= 3'b111;  
registros[2432]= 3'b100;  
registros[2433]= 3'b100;  
registros[2434]= 3'b100;  
registros[2435]= 3'b100;  
registros[2436]= 3'b100;  
registros[2437]= 3'b100;  
registros[2438]= 3'b100;  
registros[2439]= 3'b100;  
registros[2440]= 3'b100;  
registros[2441]= 3'b100;  
registros[2442]= 3'b100;  
registros[2443]= 3'b100;  
registros[2444]= 3'b100;  
registros[2445]= 3'b100;  
registros[2446]= 3'b100;  
registros[2447]= 3'b100;  
registros[2448]= 3'b100;  
registros[2449]= 3'b100;  
registros[2450]= 3'b100;  
registros[2451]= 3'b100;  
registros[2452]= 3'b100;  
registros[2453]= 3'b100;  
registros[2454]= 3'b100;  
registros[2455]= 3'b100;  
registros[2456]= 3'b100;  
registros[2457]= 3'b100;  
registros[2458]= 3'b100;  
registros[2459]= 3'b100;  
registros[2460]= 3'b100;  
registros[2461]= 3'b100;  
registros[2462]= 3'b100;  
registros[2463]= 3'b100;  
registros[2464]= 3'b100;  
registros[2465]= 3'b100;  
registros[2466]= 3'b100;  
registros[2467]= 3'b100;  
registros[2468]= 3'b100;  
registros[2469]= 3'b100;  
registros[2470]= 3'b100;  
registros[2471]= 3'b100;  
registros[2472]= 3'b100;  
registros[2473]= 3'b100;  
registros[2474]= 3'b100;  
registros[2475]= 3'b000;  
registros[2476]= 3'b100;  
registros[2477]= 3'b100;  
registros[2478]= 3'b100;  
registros[2479]= 3'b100;  
registros[2480]= 3'b100;  
registros[2481]= 3'b100;  
registros[2482]= 3'b100;  
registros[2483]= 3'b000;  
registros[2484]= 3'b000;  
registros[2485]= 3'b000;  
registros[2486]= 3'b000;  
registros[2487]= 3'b000;  
registros[2488]= 3'b000;  
registros[2489]= 3'b000;  
registros[2490]= 3'b000;  
registros[2491]= 3'b000;  
registros[2492]= 3'b000;  
registros[2493]= 3'b000;  
registros[2494]= 3'b000;  
registros[2495]= 3'b111;  
registros[2496]= 3'b000;  
registros[2497]= 3'b100;  
registros[2498]= 3'b100;  
registros[2499]= 3'b100;  
registros[2500]= 3'b100;  
registros[2501]= 3'b100;  
registros[2502]= 3'b100;  
registros[2503]= 3'b100;  
registros[2504]= 3'b110;  
registros[2505]= 3'b110;  
registros[2506]= 3'b110;  
registros[2507]= 3'b100;  
registros[2508]= 3'b100;  
registros[2509]= 3'b100;  
registros[2510]= 3'b100;  
registros[2511]= 3'b100;  
registros[2512]= 3'b100;  
registros[2513]= 3'b100;  
registros[2514]= 3'b100;  
registros[2515]= 3'b100;  
registros[2516]= 3'b100;  
registros[2517]= 3'b100;  
registros[2518]= 3'b100;  
registros[2519]= 3'b100;  
registros[2520]= 3'b100;  
registros[2521]= 3'b100;  
registros[2522]= 3'b100;  
registros[2523]= 3'b100;  
registros[2524]= 3'b100;  
registros[2525]= 3'b100;  
registros[2526]= 3'b100;  
registros[2527]= 3'b100;  
registros[2528]= 3'b100;  
registros[2529]= 3'b100;  
registros[2530]= 3'b100;  
registros[2531]= 3'b100;  
registros[2532]= 3'b100;  
registros[2533]= 3'b100;  
registros[2534]= 3'b100;  
registros[2535]= 3'b100;  
registros[2536]= 3'b100;  
registros[2537]= 3'b100;  
registros[2538]= 3'b100;  
registros[2539]= 3'b100;  
registros[2540]= 3'b100;  
registros[2541]= 3'b100;  
registros[2542]= 3'b100;  
registros[2543]= 3'b100;  
registros[2544]= 3'b100;  
registros[2545]= 3'b100;  
registros[2546]= 3'b000;  
registros[2547]= 3'b000;  
registros[2548]= 3'b000;  
registros[2549]= 3'b000;  
registros[2550]= 3'b000;  
registros[2551]= 3'b000;  
registros[2552]= 3'b000;  
registros[2553]= 3'b000;  
registros[2554]= 3'b000;  
registros[2555]= 3'b000;  
registros[2556]= 3'b000;  
registros[2557]= 3'b000;  
registros[2558]= 3'b000;  
registros[2559]= 3'b111;  
registros[2560]= 3'b111;  
registros[2561]= 3'b000;  
registros[2562]= 3'b100;  
registros[2563]= 3'b100;  
registros[2564]= 3'b100;  
registros[2565]= 3'b100;  
registros[2566]= 3'b100;  
registros[2567]= 3'b100;  
registros[2568]= 3'b110;  
registros[2569]= 3'b110;  
registros[2570]= 3'b110;  
registros[2571]= 3'b110;  
registros[2572]= 3'b110;  
registros[2573]= 3'b100;  
registros[2574]= 3'b100;  
registros[2575]= 3'b100;  
registros[2576]= 3'b100;  
registros[2577]= 3'b110;  
registros[2578]= 3'b100;  
registros[2579]= 3'b100;  
registros[2580]= 3'b100;  
registros[2581]= 3'b100;  
registros[2582]= 3'b100;  
registros[2583]= 3'b100;  
registros[2584]= 3'b100;  
registros[2585]= 3'b100;  
registros[2586]= 3'b100;  
registros[2587]= 3'b100;  
registros[2588]= 3'b100;  
registros[2589]= 3'b100;  
registros[2590]= 3'b100;  
registros[2591]= 3'b100;  
registros[2592]= 3'b100;  
registros[2593]= 3'b100;  
registros[2594]= 3'b100;  
registros[2595]= 3'b100;  
registros[2596]= 3'b100;  
registros[2597]= 3'b100;  
registros[2598]= 3'b100;  
registros[2599]= 3'b100;  
registros[2600]= 3'b100;  
registros[2601]= 3'b100;  
registros[2602]= 3'b100;  
registros[2603]= 3'b100;  
registros[2604]= 3'b100;  
registros[2605]= 3'b100;  
registros[2606]= 3'b100;  
registros[2607]= 3'b000;  
registros[2608]= 3'b100;  
registros[2609]= 3'b100;  
registros[2610]= 3'b000;  
registros[2611]= 3'b000;  
registros[2612]= 3'b000;  
registros[2613]= 3'b000;  
registros[2614]= 3'b000;  
registros[2615]= 3'b000;  
registros[2616]= 3'b000;  
registros[2617]= 3'b000;  
registros[2618]= 3'b000;  
registros[2619]= 3'b000;  
registros[2620]= 3'b000;  
registros[2621]= 3'b000;  
registros[2622]= 3'b000;  
registros[2623]= 3'b111;  
registros[2624]= 3'b111;  
registros[2625]= 3'b111;  
registros[2626]= 3'b100;  
registros[2627]= 3'b100;  
registros[2628]= 3'b100;  
registros[2629]= 3'b100;  
registros[2630]= 3'b100;  
registros[2631]= 3'b100;  
registros[2632]= 3'b100;  
registros[2633]= 3'b100;  
registros[2634]= 3'b100;  
registros[2635]= 3'b110;  
registros[2636]= 3'b110;  
registros[2637]= 3'b110;  
registros[2638]= 3'b100;  
registros[2639]= 3'b110;  
registros[2640]= 3'b110;  
registros[2641]= 3'b110;  
registros[2642]= 3'b100;  
registros[2643]= 3'b100;  
registros[2644]= 3'b110;  
registros[2645]= 3'b100;  
registros[2646]= 3'b100;  
registros[2647]= 3'b110;  
registros[2648]= 3'b100;  
registros[2649]= 3'b100;  
registros[2650]= 3'b100;  
registros[2651]= 3'b100;  
registros[2652]= 3'b100;  
registros[2653]= 3'b100;  
registros[2654]= 3'b100;  
registros[2655]= 3'b100;  
registros[2656]= 3'b100;  
registros[2657]= 3'b100;  
registros[2658]= 3'b100;  
registros[2659]= 3'b100;  
registros[2660]= 3'b100;  
registros[2661]= 3'b100;  
registros[2662]= 3'b100;  
registros[2663]= 3'b100;  
registros[2664]= 3'b100;  
registros[2665]= 3'b100;  
registros[2666]= 3'b100;  
registros[2667]= 3'b100;  
registros[2668]= 3'b100;  
registros[2669]= 3'b100;  
registros[2670]= 3'b100;  
registros[2671]= 3'b100;  
registros[2672]= 3'b100;  
registros[2673]= 3'b100;  
registros[2674]= 3'b100;  
registros[2675]= 3'b000;  
registros[2676]= 3'b000;  
registros[2677]= 3'b000;  
registros[2678]= 3'b100;  
registros[2679]= 3'b000;  
registros[2680]= 3'b000;  
registros[2681]= 3'b000;  
registros[2682]= 3'b000;  
registros[2683]= 3'b000;  
registros[2684]= 3'b000;  
registros[2685]= 3'b000;  
registros[2686]= 3'b000;  
registros[2687]= 3'b111;  
registros[2688]= 3'b111;  
registros[2689]= 3'b111;  
registros[2690]= 3'b000;  
registros[2691]= 3'b000;  
registros[2692]= 3'b000;  
registros[2693]= 3'b100;  
registros[2694]= 3'b100;  
registros[2695]= 3'b100;  
registros[2696]= 3'b100;  
registros[2697]= 3'b100;  
registros[2698]= 3'b100;  
registros[2699]= 3'b100;  
registros[2700]= 3'b100;  
registros[2701]= 3'b110;  
registros[2702]= 3'b100;  
registros[2703]= 3'b110;  
registros[2704]= 3'b110;  
registros[2705]= 3'b100;  
registros[2706]= 3'b100;  
registros[2707]= 3'b100;  
registros[2708]= 3'b100;  
registros[2709]= 3'b110;  
registros[2710]= 3'b110;  
registros[2711]= 3'b110;  
registros[2712]= 3'b110;  
registros[2713]= 3'b100;  
registros[2714]= 3'b100;  
registros[2715]= 3'b100;  
registros[2716]= 3'b100;  
registros[2717]= 3'b100;  
registros[2718]= 3'b100;  
registros[2719]= 3'b100;  
registros[2720]= 3'b100;  
registros[2721]= 3'b100;  
registros[2722]= 3'b100;  
registros[2723]= 3'b100;  
registros[2724]= 3'b100;  
registros[2725]= 3'b100;  
registros[2726]= 3'b100;  
registros[2727]= 3'b100;  
registros[2728]= 3'b100;  
registros[2729]= 3'b100;  
registros[2730]= 3'b100;  
registros[2731]= 3'b100;  
registros[2732]= 3'b100;  
registros[2733]= 3'b100;  
registros[2734]= 3'b100;  
registros[2735]= 3'b100;  
registros[2736]= 3'b100;  
registros[2737]= 3'b100;  
registros[2738]= 3'b100;  
registros[2739]= 3'b100;  
registros[2740]= 3'b100;  
registros[2741]= 3'b000;  
registros[2742]= 3'b000;  
registros[2743]= 3'b000;  
registros[2744]= 3'b000;  
registros[2745]= 3'b000;  
registros[2746]= 3'b000;  
registros[2747]= 3'b000;  
registros[2748]= 3'b000;  
registros[2749]= 3'b111;  
registros[2750]= 3'b111;  
registros[2751]= 3'b111;  
registros[2752]= 3'b111;  
registros[2753]= 3'b111;  
registros[2754]= 3'b111;  
registros[2755]= 3'b000;  
registros[2756]= 3'b000;  
registros[2757]= 3'b000;  
registros[2758]= 3'b000;  
registros[2759]= 3'b100;  
registros[2760]= 3'b100;  
registros[2761]= 3'b100;  
registros[2762]= 3'b100;  
registros[2763]= 3'b100;  
registros[2764]= 3'b100;  
registros[2765]= 3'b100;  
registros[2766]= 3'b100;  
registros[2767]= 3'b110;  
registros[2768]= 3'b100;  
registros[2769]= 3'b100;  
registros[2770]= 3'b100;  
registros[2771]= 3'b100;  
registros[2772]= 3'b100;  
registros[2773]= 3'b110;  
registros[2774]= 3'b110;  
registros[2775]= 3'b110;  
registros[2776]= 3'b110;  
registros[2777]= 3'b100;  
registros[2778]= 3'b100;  
registros[2779]= 3'b100;  
registros[2780]= 3'b100;  
registros[2781]= 3'b100;  
registros[2782]= 3'b100;  
registros[2783]= 3'b100;  
registros[2784]= 3'b100;  
registros[2785]= 3'b100;  
registros[2786]= 3'b100;  
registros[2787]= 3'b100;  
registros[2788]= 3'b100;  
registros[2789]= 3'b100;  
registros[2790]= 3'b100;  
registros[2791]= 3'b100;  
registros[2792]= 3'b100;  
registros[2793]= 3'b100;  
registros[2794]= 3'b100;  
registros[2795]= 3'b100;  
registros[2796]= 3'b100;  
registros[2797]= 3'b100;  
registros[2798]= 3'b000;  
registros[2799]= 3'b000;  
registros[2800]= 3'b100;  
registros[2801]= 3'b100;  
registros[2802]= 3'b100;  
registros[2803]= 3'b100;  
registros[2804]= 3'b100;  
registros[2805]= 3'b100;  
registros[2806]= 3'b000;  
registros[2807]= 3'b000;  
registros[2808]= 3'b000;  
registros[2809]= 3'b000;  
registros[2810]= 3'b000;  
registros[2811]= 3'b000;  
registros[2812]= 3'b111;  
registros[2813]= 3'b111;  
registros[2814]= 3'b111;  
registros[2815]= 3'b111;  
registros[2816]= 3'b111;  
registros[2817]= 3'b111;  
registros[2818]= 3'b111;  
registros[2819]= 3'b111;  
registros[2820]= 3'b000;  
registros[2821]= 3'b000;  
registros[2822]= 3'b000;  
registros[2823]= 3'b100;  
registros[2824]= 3'b100;  
registros[2825]= 3'b100;  
registros[2826]= 3'b100;  
registros[2827]= 3'b100;  
registros[2828]= 3'b100;  
registros[2829]= 3'b100;  
registros[2830]= 3'b100;  
registros[2831]= 3'b110;  
registros[2832]= 3'b110;  
registros[2833]= 3'b110;  
registros[2834]= 3'b110;  
registros[2835]= 3'b110;  
registros[2836]= 3'b110;  
registros[2837]= 3'b110;  
registros[2838]= 3'b110;  
registros[2839]= 3'b110;  
registros[2840]= 3'b110;  
registros[2841]= 3'b100;  
registros[2842]= 3'b100;  
registros[2843]= 3'b100;  
registros[2844]= 3'b100;  
registros[2845]= 3'b100;  
registros[2846]= 3'b100;  
registros[2847]= 3'b100;  
registros[2848]= 3'b100;  
registros[2849]= 3'b100;  
registros[2850]= 3'b100;  
registros[2851]= 3'b100;  
registros[2852]= 3'b100;  
registros[2853]= 3'b100;  
registros[2854]= 3'b100;  
registros[2855]= 3'b100;  
registros[2856]= 3'b100;  
registros[2857]= 3'b100;  
registros[2858]= 3'b100;  
registros[2859]= 3'b100;  
registros[2860]= 3'b100;  
registros[2861]= 3'b100;  
registros[2862]= 3'b000;  
registros[2863]= 3'b100;  
registros[2864]= 3'b100;  
registros[2865]= 3'b100;  
registros[2866]= 3'b100;  
registros[2867]= 3'b100;  
registros[2868]= 3'b100;  
registros[2869]= 3'b000;  
registros[2870]= 3'b000;  
registros[2871]= 3'b000;  
registros[2872]= 3'b000;  
registros[2873]= 3'b000;  
registros[2874]= 3'b000;  
registros[2875]= 3'b111;  
registros[2876]= 3'b111;  
registros[2877]= 3'b111;  
registros[2878]= 3'b111;  
registros[2879]= 3'b111;  
registros[2880]= 3'b111;  
registros[2881]= 3'b111;  
registros[2882]= 3'b111;  
registros[2883]= 3'b111;  
registros[2884]= 3'b111;  
registros[2885]= 3'b000;  
registros[2886]= 3'b100;  
registros[2887]= 3'b100;  
registros[2888]= 3'b100;  
registros[2889]= 3'b100;  
registros[2890]= 3'b100;  
registros[2891]= 3'b100;  
registros[2892]= 3'b100;  
registros[2893]= 3'b100;  
registros[2894]= 3'b100;  
registros[2895]= 3'b110;  
registros[2896]= 3'b110;  
registros[2897]= 3'b110;  
registros[2898]= 3'b110;  
registros[2899]= 3'b110;  
registros[2900]= 3'b110;  
registros[2901]= 3'b110;  
registros[2902]= 3'b110;  
registros[2903]= 3'b110;  
registros[2904]= 3'b100;  
registros[2905]= 3'b100;  
registros[2906]= 3'b100;  
registros[2907]= 3'b100;  
registros[2908]= 3'b100;  
registros[2909]= 3'b100;  
registros[2910]= 3'b100;  
registros[2911]= 3'b100;  
registros[2912]= 3'b100;  
registros[2913]= 3'b100;  
registros[2914]= 3'b100;  
registros[2915]= 3'b100;  
registros[2916]= 3'b100;  
registros[2917]= 3'b100;  
registros[2918]= 3'b100;  
registros[2919]= 3'b100;  
registros[2920]= 3'b100;  
registros[2921]= 3'b100;  
registros[2922]= 3'b100;  
registros[2923]= 3'b100;  
registros[2924]= 3'b100;  
registros[2925]= 3'b100;  
registros[2926]= 3'b100;  
registros[2927]= 3'b100;  
registros[2928]= 3'b100;  
registros[2929]= 3'b100;  
registros[2930]= 3'b100;  
registros[2931]= 3'b100;  
registros[2932]= 3'b100;  
registros[2933]= 3'b000;  
registros[2934]= 3'b000;  
registros[2935]= 3'b000;  
registros[2936]= 3'b000;  
registros[2937]= 3'b000;  
registros[2938]= 3'b111;  
registros[2939]= 3'b111;  
registros[2940]= 3'b111;  
registros[2941]= 3'b111;  
registros[2942]= 3'b111;  
registros[2943]= 3'b111;  
registros[2944]= 3'b111;  
registros[2945]= 3'b111;  
registros[2946]= 3'b111;  
registros[2947]= 3'b111;  
registros[2948]= 3'b111;  
registros[2949]= 3'b000;  
registros[2950]= 3'b100;  
registros[2951]= 3'b100;  
registros[2952]= 3'b100;  
registros[2953]= 3'b100;  
registros[2954]= 3'b100;  
registros[2955]= 3'b100;  
registros[2956]= 3'b100;  
registros[2957]= 3'b100;  
registros[2958]= 3'b100;  
registros[2959]= 3'b100;  
registros[2960]= 3'b110;  
registros[2961]= 3'b110;  
registros[2962]= 3'b110;  
registros[2963]= 3'b110;  
registros[2964]= 3'b110;  
registros[2965]= 3'b110;  
registros[2966]= 3'b110;  
registros[2967]= 3'b100;  
registros[2968]= 3'b100;  
registros[2969]= 3'b100;  
registros[2970]= 3'b100;  
registros[2971]= 3'b100;  
registros[2972]= 3'b100;  
registros[2973]= 3'b100;  
registros[2974]= 3'b100;  
registros[2975]= 3'b100;  
registros[2976]= 3'b100;  
registros[2977]= 3'b100;  
registros[2978]= 3'b100;  
registros[2979]= 3'b100;  
registros[2980]= 3'b100;  
registros[2981]= 3'b100;  
registros[2982]= 3'b100;  
registros[2983]= 3'b100;  
registros[2984]= 3'b100;  
registros[2985]= 3'b100;  
registros[2986]= 3'b100;  
registros[2987]= 3'b100;  
registros[2988]= 3'b100;  
registros[2989]= 3'b100;  
registros[2990]= 3'b100;  
registros[2991]= 3'b100;  
registros[2992]= 3'b100;  
registros[2993]= 3'b100;  
registros[2994]= 3'b100;  
registros[2995]= 3'b100;  
registros[2996]= 3'b000;  
registros[2997]= 3'b000;  
registros[2998]= 3'b000;  
registros[2999]= 3'b000;  
registros[3000]= 3'b000;  
registros[3001]= 3'b000;  
registros[3002]= 3'b111;  
registros[3003]= 3'b111;  
registros[3004]= 3'b111;  
registros[3005]= 3'b111;  
registros[3006]= 3'b111;  
registros[3007]= 3'b111;  
registros[3008]= 3'b111;  
registros[3009]= 3'b111;  
registros[3010]= 3'b111;  
registros[3011]= 3'b111;  
registros[3012]= 3'b111;  
registros[3013]= 3'b111;  
registros[3014]= 3'b000;  
registros[3015]= 3'b100;  
registros[3016]= 3'b100;  
registros[3017]= 3'b100;  
registros[3018]= 3'b100;  
registros[3019]= 3'b100;  
registros[3020]= 3'b100;  
registros[3021]= 3'b100;  
registros[3022]= 3'b100;  
registros[3023]= 3'b100;  
registros[3024]= 3'b110;  
registros[3025]= 3'b110;  
registros[3026]= 3'b110;  
registros[3027]= 3'b110;  
registros[3028]= 3'b110;  
registros[3029]= 3'b110;  
registros[3030]= 3'b110;  
registros[3031]= 3'b100;  
registros[3032]= 3'b100;  
registros[3033]= 3'b100;  
registros[3034]= 3'b100;  
registros[3035]= 3'b100;  
registros[3036]= 3'b100;  
registros[3037]= 3'b100;  
registros[3038]= 3'b100;  
registros[3039]= 3'b100;  
registros[3040]= 3'b100;  
registros[3041]= 3'b100;  
registros[3042]= 3'b000;  
registros[3043]= 3'b100;  
registros[3044]= 3'b100;  
registros[3045]= 3'b100;  
registros[3046]= 3'b100;  
registros[3047]= 3'b100;  
registros[3048]= 3'b100;  
registros[3049]= 3'b100;  
registros[3050]= 3'b100;  
registros[3051]= 3'b100;  
registros[3052]= 3'b100;  
registros[3053]= 3'b100;  
registros[3054]= 3'b100;  
registros[3055]= 3'b100;  
registros[3056]= 3'b100;  
registros[3057]= 3'b100;  
registros[3058]= 3'b100;  
registros[3059]= 3'b100;  
registros[3060]= 3'b000;  
registros[3061]= 3'b000;  
registros[3062]= 3'b000;  
registros[3063]= 3'b000;  
registros[3064]= 3'b000;  
registros[3065]= 3'b000;  
registros[3066]= 3'b111;  
registros[3067]= 3'b111;  
registros[3068]= 3'b111;  
registros[3069]= 3'b111;  
registros[3070]= 3'b111;  
registros[3071]= 3'b111;  
registros[3072]= 3'b111;  
registros[3073]= 3'b111;  
registros[3074]= 3'b111;  
registros[3075]= 3'b111;  
registros[3076]= 3'b111;  
registros[3077]= 3'b111;  
registros[3078]= 3'b111;  
registros[3079]= 3'b000;  
registros[3080]= 3'b100;  
registros[3081]= 3'b100;  
registros[3082]= 3'b100;  
registros[3083]= 3'b100;  
registros[3084]= 3'b100;  
registros[3085]= 3'b100;  
registros[3086]= 3'b100;  
registros[3087]= 3'b100;  
registros[3088]= 3'b100;  
registros[3089]= 3'b110;  
registros[3090]= 3'b110;  
registros[3091]= 3'b110;  
registros[3092]= 3'b110;  
registros[3093]= 3'b110;  
registros[3094]= 3'b110;  
registros[3095]= 3'b100;  
registros[3096]= 3'b100;  
registros[3097]= 3'b100;  
registros[3098]= 3'b100;  
registros[3099]= 3'b100;  
registros[3100]= 3'b100;  
registros[3101]= 3'b100;  
registros[3102]= 3'b100;  
registros[3103]= 3'b100;  
registros[3104]= 3'b100;  
registros[3105]= 3'b100;  
registros[3106]= 3'b000;  
registros[3107]= 3'b100;  
registros[3108]= 3'b100;  
registros[3109]= 3'b100;  
registros[3110]= 3'b100;  
registros[3111]= 3'b100;  
registros[3112]= 3'b100;  
registros[3113]= 3'b100;  
registros[3114]= 3'b100;  
registros[3115]= 3'b100;  
registros[3116]= 3'b100;  
registros[3117]= 3'b100;  
registros[3118]= 3'b100;  
registros[3119]= 3'b100;  
registros[3120]= 3'b100;  
registros[3121]= 3'b100;  
registros[3122]= 3'b100;  
registros[3123]= 3'b100;  
registros[3124]= 3'b000;  
registros[3125]= 3'b000;  
registros[3126]= 3'b000;  
registros[3127]= 3'b000;  
registros[3128]= 3'b000;  
registros[3129]= 3'b000;  
registros[3130]= 3'b111;  
registros[3131]= 3'b111;  
registros[3132]= 3'b111;  
registros[3133]= 3'b111;  
registros[3134]= 3'b111;  
registros[3135]= 3'b111;  
registros[3136]= 3'b111;  
registros[3137]= 3'b111;  
registros[3138]= 3'b111;  
registros[3139]= 3'b111;  
registros[3140]= 3'b111;  
registros[3141]= 3'b111;  
registros[3142]= 3'b111;  
registros[3143]= 3'b000;  
registros[3144]= 3'b000;  
registros[3145]= 3'b100;  
registros[3146]= 3'b000;  
registros[3147]= 3'b000;  
registros[3148]= 3'b100;  
registros[3149]= 3'b100;  
registros[3150]= 3'b100;  
registros[3151]= 3'b100;  
registros[3152]= 3'b100;  
registros[3153]= 3'b100;  
registros[3154]= 3'b110;  
registros[3155]= 3'b110;  
registros[3156]= 3'b110;  
registros[3157]= 3'b110;  
registros[3158]= 3'b100;  
registros[3159]= 3'b100;  
registros[3160]= 3'b100;  
registros[3161]= 3'b100;  
registros[3162]= 3'b100;  
registros[3163]= 3'b100;  
registros[3164]= 3'b100;  
registros[3165]= 3'b100;  
registros[3166]= 3'b100;  
registros[3167]= 3'b100;  
registros[3168]= 3'b100;  
registros[3169]= 3'b000;  
registros[3170]= 3'b000;  
registros[3171]= 3'b000;  
registros[3172]= 3'b000;  
registros[3173]= 3'b000;  
registros[3174]= 3'b000;  
registros[3175]= 3'b000;  
registros[3176]= 3'b000;  
registros[3177]= 3'b000;  
registros[3178]= 3'b000;  
registros[3179]= 3'b100;  
registros[3180]= 3'b100;  
registros[3181]= 3'b100;  
registros[3182]= 3'b100;  
registros[3183]= 3'b100;  
registros[3184]= 3'b100;  
registros[3185]= 3'b100;  
registros[3186]= 3'b100;  
registros[3187]= 3'b100;  
registros[3188]= 3'b000;  
registros[3189]= 3'b000;  
registros[3190]= 3'b000;  
registros[3191]= 3'b000;  
registros[3192]= 3'b000;  
registros[3193]= 3'b111;  
registros[3194]= 3'b111;  
registros[3195]= 3'b111;  
registros[3196]= 3'b111;  
registros[3197]= 3'b111;  
registros[3198]= 3'b111;  
registros[3199]= 3'b111;  
registros[3200]= 3'b111;  
registros[3201]= 3'b111;  
registros[3202]= 3'b111;  
registros[3203]= 3'b111;  
registros[3204]= 3'b111;  
registros[3205]= 3'b111;  
registros[3206]= 3'b111;  
registros[3207]= 3'b111;  
registros[3208]= 3'b000;  
registros[3209]= 3'b000;  
registros[3210]= 3'b000;  
registros[3211]= 3'b000;  
registros[3212]= 3'b100;  
registros[3213]= 3'b100;  
registros[3214]= 3'b100;  
registros[3215]= 3'b100;  
registros[3216]= 3'b100;  
registros[3217]= 3'b100;  
registros[3218]= 3'b100;  
registros[3219]= 3'b100;  
registros[3220]= 3'b100;  
registros[3221]= 3'b100;  
registros[3222]= 3'b100;  
registros[3223]= 3'b100;  
registros[3224]= 3'b100;  
registros[3225]= 3'b100;  
registros[3226]= 3'b100;  
registros[3227]= 3'b100;  
registros[3228]= 3'b100;  
registros[3229]= 3'b100;  
registros[3230]= 3'b100;  
registros[3231]= 3'b100;  
registros[3232]= 3'b100;  
registros[3233]= 3'b000;  
registros[3234]= 3'b100;  
registros[3235]= 3'b000;  
registros[3236]= 3'b000;  
registros[3237]= 3'b000;  
registros[3238]= 3'b000;  
registros[3239]= 3'b000;  
registros[3240]= 3'b000;  
registros[3241]= 3'b000;  
registros[3242]= 3'b000;  
registros[3243]= 3'b000;  
registros[3244]= 3'b100;  
registros[3245]= 3'b100;  
registros[3246]= 3'b100;  
registros[3247]= 3'b100;  
registros[3248]= 3'b100;  
registros[3249]= 3'b100;  
registros[3250]= 3'b000;  
registros[3251]= 3'b000;  
registros[3252]= 3'b000;  
registros[3253]= 3'b000;  
registros[3254]= 3'b000;  
registros[3255]= 3'b000;  
registros[3256]= 3'b000;  
registros[3257]= 3'b111;  
registros[3258]= 3'b111;  
registros[3259]= 3'b111;  
registros[3260]= 3'b111;  
registros[3261]= 3'b111;  
registros[3262]= 3'b111;  
registros[3263]= 3'b111;  
registros[3264]= 3'b111;  
registros[3265]= 3'b111;  
registros[3266]= 3'b111;  
registros[3267]= 3'b111;  
registros[3268]= 3'b111;  
registros[3269]= 3'b111;  
registros[3270]= 3'b111;  
registros[3271]= 3'b111;  
registros[3272]= 3'b000;  
registros[3273]= 3'b000;  
registros[3274]= 3'b000;  
registros[3275]= 3'b000;  
registros[3276]= 3'b100;  
registros[3277]= 3'b100;  
registros[3278]= 3'b100;  
registros[3279]= 3'b100;  
registros[3280]= 3'b100;  
registros[3281]= 3'b100;  
registros[3282]= 3'b100;  
registros[3283]= 3'b100;  
registros[3284]= 3'b100;  
registros[3285]= 3'b100;  
registros[3286]= 3'b100;  
registros[3287]= 3'b100;  
registros[3288]= 3'b100;  
registros[3289]= 3'b100;  
registros[3290]= 3'b100;  
registros[3291]= 3'b100;  
registros[3292]= 3'b100;  
registros[3293]= 3'b100;  
registros[3294]= 3'b100;  
registros[3295]= 3'b100;  
registros[3296]= 3'b100;  
registros[3297]= 3'b100;  
registros[3298]= 3'b100;  
registros[3299]= 3'b100;  
registros[3300]= 3'b000;  
registros[3301]= 3'b000;  
registros[3302]= 3'b000;  
registros[3303]= 3'b000;  
registros[3304]= 3'b000;  
registros[3305]= 3'b000;  
registros[3306]= 3'b000;  
registros[3307]= 3'b000;  
registros[3308]= 3'b000;  
registros[3309]= 3'b000;  
registros[3310]= 3'b100;  
registros[3311]= 3'b100;  
registros[3312]= 3'b100;  
registros[3313]= 3'b100;  
registros[3314]= 3'b100;  
registros[3315]= 3'b000;  
registros[3316]= 3'b000;  
registros[3317]= 3'b000;  
registros[3318]= 3'b000;  
registros[3319]= 3'b000;  
registros[3320]= 3'b111;  
registros[3321]= 3'b111;  
registros[3322]= 3'b111;  
registros[3323]= 3'b111;  
registros[3324]= 3'b111;  
registros[3325]= 3'b111;  
registros[3326]= 3'b111;  
registros[3327]= 3'b111;  
registros[3328]= 3'b111;  
registros[3329]= 3'b111;  
registros[3330]= 3'b111;  
registros[3331]= 3'b111;  
registros[3332]= 3'b111;  
registros[3333]= 3'b111;  
registros[3334]= 3'b111;  
registros[3335]= 3'b111;  
registros[3336]= 3'b000;  
registros[3337]= 3'b000;  
registros[3338]= 3'b000;  
registros[3339]= 3'b100;  
registros[3340]= 3'b100;  
registros[3341]= 3'b100;  
registros[3342]= 3'b100;  
registros[3343]= 3'b100;  
registros[3344]= 3'b100;  
registros[3345]= 3'b100;  
registros[3346]= 3'b100;  
registros[3347]= 3'b100;  
registros[3348]= 3'b100;  
registros[3349]= 3'b100;  
registros[3350]= 3'b100;  
registros[3351]= 3'b100;  
registros[3352]= 3'b100;  
registros[3353]= 3'b100;  
registros[3354]= 3'b100;  
registros[3355]= 3'b100;  
registros[3356]= 3'b100;  
registros[3357]= 3'b100;  
registros[3358]= 3'b100;  
registros[3359]= 3'b100;  
registros[3360]= 3'b100;  
registros[3361]= 3'b100;  
registros[3362]= 3'b100;  
registros[3363]= 3'b000;  
registros[3364]= 3'b000;  
registros[3365]= 3'b000;  
registros[3366]= 3'b000;  
registros[3367]= 3'b000;  
registros[3368]= 3'b000;  
registros[3369]= 3'b000;  
registros[3370]= 3'b000;  
registros[3371]= 3'b000;  
registros[3372]= 3'b000;  
registros[3373]= 3'b000;  
registros[3374]= 3'b000;  
registros[3375]= 3'b100;  
registros[3376]= 3'b100;  
registros[3377]= 3'b100;  
registros[3378]= 3'b100;  
registros[3379]= 3'b000;  
registros[3380]= 3'b000;  
registros[3381]= 3'b000;  
registros[3382]= 3'b000;  
registros[3383]= 3'b111;  
registros[3384]= 3'b111;  
registros[3385]= 3'b111;  
registros[3386]= 3'b111;  
registros[3387]= 3'b111;  
registros[3388]= 3'b111;  
registros[3389]= 3'b111;  
registros[3390]= 3'b111;  
registros[3391]= 3'b111;  
registros[3392]= 3'b111;  
registros[3393]= 3'b111;  
registros[3394]= 3'b111;  
registros[3395]= 3'b111;  
registros[3396]= 3'b111;  
registros[3397]= 3'b111;  
registros[3398]= 3'b111;  
registros[3399]= 3'b111;  
registros[3400]= 3'b000;  
registros[3401]= 3'b000;  
registros[3402]= 3'b100;  
registros[3403]= 3'b100;  
registros[3404]= 3'b100;  
registros[3405]= 3'b100;  
registros[3406]= 3'b100;  
registros[3407]= 3'b100;  
registros[3408]= 3'b100;  
registros[3409]= 3'b100;  
registros[3410]= 3'b100;  
registros[3411]= 3'b100;  
registros[3412]= 3'b100;  
registros[3413]= 3'b100;  
registros[3414]= 3'b100;  
registros[3415]= 3'b100;  
registros[3416]= 3'b100;  
registros[3417]= 3'b100;  
registros[3418]= 3'b100;  
registros[3419]= 3'b100;  
registros[3420]= 3'b100;  
registros[3421]= 3'b100;  
registros[3422]= 3'b100;  
registros[3423]= 3'b100;  
registros[3424]= 3'b100;  
registros[3425]= 3'b100;  
registros[3426]= 3'b100;  
registros[3427]= 3'b000;  
registros[3428]= 3'b000;  
registros[3429]= 3'b000;  
registros[3430]= 3'b000;  
registros[3431]= 3'b000;  
registros[3432]= 3'b000;  
registros[3433]= 3'b000;  
registros[3434]= 3'b000;  
registros[3435]= 3'b000;  
registros[3436]= 3'b000;  
registros[3437]= 3'b000;  
registros[3438]= 3'b000;  
registros[3439]= 3'b000;  
registros[3440]= 3'b000;  
registros[3441]= 3'b100;  
registros[3442]= 3'b100;  
registros[3443]= 3'b000;  
registros[3444]= 3'b000;  
registros[3445]= 3'b111;  
registros[3446]= 3'b111;  
registros[3447]= 3'b111;  
registros[3448]= 3'b111;  
registros[3449]= 3'b111;  
registros[3450]= 3'b111;  
registros[3451]= 3'b111;  
registros[3452]= 3'b111;  
registros[3453]= 3'b111;  
registros[3454]= 3'b111;  
registros[3455]= 3'b111;  
registros[3456]= 3'b111;  
registros[3457]= 3'b111;  
registros[3458]= 3'b111;  
registros[3459]= 3'b111;  
registros[3460]= 3'b111;  
registros[3461]= 3'b111;  
registros[3462]= 3'b111;  
registros[3463]= 3'b111;  
registros[3464]= 3'b111;  
registros[3465]= 3'b000;  
registros[3466]= 3'b000;  
registros[3467]= 3'b100;  
registros[3468]= 3'b100;  
registros[3469]= 3'b100;  
registros[3470]= 3'b100;  
registros[3471]= 3'b100;  
registros[3472]= 3'b100;  
registros[3473]= 3'b100;  
registros[3474]= 3'b100;  
registros[3475]= 3'b100;  
registros[3476]= 3'b100;  
registros[3477]= 3'b100;  
registros[3478]= 3'b100;  
registros[3479]= 3'b100;  
registros[3480]= 3'b100;  
registros[3481]= 3'b100;  
registros[3482]= 3'b100;  
registros[3483]= 3'b100;  
registros[3484]= 3'b100;  
registros[3485]= 3'b100;  
registros[3486]= 3'b100;  
registros[3487]= 3'b100;  
registros[3488]= 3'b100;  
registros[3489]= 3'b100;  
registros[3490]= 3'b100;  
registros[3491]= 3'b000;  
registros[3492]= 3'b000;  
registros[3493]= 3'b000;  
registros[3494]= 3'b000;  
registros[3495]= 3'b000;  
registros[3496]= 3'b000;  
registros[3497]= 3'b000;  
registros[3498]= 3'b000;  
registros[3499]= 3'b000;  
registros[3500]= 3'b000;  
registros[3501]= 3'b000;  
registros[3502]= 3'b000;  
registros[3503]= 3'b000;  
registros[3504]= 3'b000;  
registros[3505]= 3'b100;  
registros[3506]= 3'b000;  
registros[3507]= 3'b000;  
registros[3508]= 3'b111;  
registros[3509]= 3'b111;  
registros[3510]= 3'b111;  
registros[3511]= 3'b111;  
registros[3512]= 3'b111;  
registros[3513]= 3'b111;  
registros[3514]= 3'b111;  
registros[3515]= 3'b111;  
registros[3516]= 3'b111;  
registros[3517]= 3'b111;  
registros[3518]= 3'b111;  
registros[3519]= 3'b111;  
registros[3520]= 3'b111;  
registros[3521]= 3'b111;  
registros[3522]= 3'b111;  
registros[3523]= 3'b111;  
registros[3524]= 3'b111;  
registros[3525]= 3'b111;  
registros[3526]= 3'b111;  
registros[3527]= 3'b111;  
registros[3528]= 3'b111;  
registros[3529]= 3'b000;  
registros[3530]= 3'b000;  
registros[3531]= 3'b000;  
registros[3532]= 3'b000;  
registros[3533]= 3'b100;  
registros[3534]= 3'b100;  
registros[3535]= 3'b100;  
registros[3536]= 3'b100;  
registros[3537]= 3'b100;  
registros[3538]= 3'b100;  
registros[3539]= 3'b100;  
registros[3540]= 3'b100;  
registros[3541]= 3'b100;  
registros[3542]= 3'b100;  
registros[3543]= 3'b100;  
registros[3544]= 3'b100;  
registros[3545]= 3'b100;  
registros[3546]= 3'b100;  
registros[3547]= 3'b100;  
registros[3548]= 3'b100;  
registros[3549]= 3'b100;  
registros[3550]= 3'b100;  
registros[3551]= 3'b100;  
registros[3552]= 3'b100;  
registros[3553]= 3'b100;  
registros[3554]= 3'b100;  
registros[3555]= 3'b100;  
registros[3556]= 3'b000;  
registros[3557]= 3'b000;  
registros[3558]= 3'b000;  
registros[3559]= 3'b000;  
registros[3560]= 3'b000;  
registros[3561]= 3'b000;  
registros[3562]= 3'b000;  
registros[3563]= 3'b000;  
registros[3564]= 3'b000;  
registros[3565]= 3'b000;  
registros[3566]= 3'b000;  
registros[3567]= 3'b000;  
registros[3568]= 3'b000;  
registros[3569]= 3'b000;  
registros[3570]= 3'b000;  
registros[3571]= 3'b111;  
registros[3572]= 3'b111;  
registros[3573]= 3'b111;  
registros[3574]= 3'b111;  
registros[3575]= 3'b111;  
registros[3576]= 3'b111;  
registros[3577]= 3'b111;  
registros[3578]= 3'b111;  
registros[3579]= 3'b111;  
registros[3580]= 3'b111;  
registros[3581]= 3'b111;  
registros[3582]= 3'b111;  
registros[3583]= 3'b111;  
registros[3584]= 3'b111;  
registros[3585]= 3'b111;  
registros[3586]= 3'b111;  
registros[3587]= 3'b111;  
registros[3588]= 3'b111;  
registros[3589]= 3'b111;  
registros[3590]= 3'b111;  
registros[3591]= 3'b111;  
registros[3592]= 3'b111;  
registros[3593]= 3'b000;  
registros[3594]= 3'b000;  
registros[3595]= 3'b000;  
registros[3596]= 3'b000;  
registros[3597]= 3'b100;  
registros[3598]= 3'b100;  
registros[3599]= 3'b100;  
registros[3600]= 3'b100;  
registros[3601]= 3'b100;  
registros[3602]= 3'b100;  
registros[3603]= 3'b100;  
registros[3604]= 3'b100;  
registros[3605]= 3'b100;  
registros[3606]= 3'b100;  
registros[3607]= 3'b100;  
registros[3608]= 3'b100;  
registros[3609]= 3'b100;  
registros[3610]= 3'b100;  
registros[3611]= 3'b100;  
registros[3612]= 3'b100;  
registros[3613]= 3'b100;  
registros[3614]= 3'b100;  
registros[3615]= 3'b100;  
registros[3616]= 3'b000;  
registros[3617]= 3'b000;  
registros[3618]= 3'b000;  
registros[3619]= 3'b000;  
registros[3620]= 3'b000;  
registros[3621]= 3'b000;  
registros[3622]= 3'b000;  
registros[3623]= 3'b000;  
registros[3624]= 3'b000;  
registros[3625]= 3'b000;  
registros[3626]= 3'b000;  
registros[3627]= 3'b000;  
registros[3628]= 3'b111;  
registros[3629]= 3'b111;  
registros[3630]= 3'b111;  
registros[3631]= 3'b111;  
registros[3632]= 3'b000;  
registros[3633]= 3'b000;  
registros[3634]= 3'b000;  
registros[3635]= 3'b111;  
registros[3636]= 3'b111;  
registros[3637]= 3'b111;  
registros[3638]= 3'b111;  
registros[3639]= 3'b111;  
registros[3640]= 3'b111;  
registros[3641]= 3'b111;  
registros[3642]= 3'b111;  
registros[3643]= 3'b111;  
registros[3644]= 3'b111;  
registros[3645]= 3'b111;  
registros[3646]= 3'b111;  
registros[3647]= 3'b111;  
registros[3648]= 3'b111;  
registros[3649]= 3'b111;  
registros[3650]= 3'b111;  
registros[3651]= 3'b111;  
registros[3652]= 3'b111;  
registros[3653]= 3'b111;  
registros[3654]= 3'b111;  
registros[3655]= 3'b111;  
registros[3656]= 3'b111;  
registros[3657]= 3'b111;  
registros[3658]= 3'b000;  
registros[3659]= 3'b000;  
registros[3660]= 3'b000;  
registros[3661]= 3'b000;  
registros[3662]= 3'b100;  
registros[3663]= 3'b100;  
registros[3664]= 3'b100;  
registros[3665]= 3'b100;  
registros[3666]= 3'b100;  
registros[3667]= 3'b000;  
registros[3668]= 3'b100;  
registros[3669]= 3'b100;  
registros[3670]= 3'b100;  
registros[3671]= 3'b100;  
registros[3672]= 3'b100;  
registros[3673]= 3'b100;  
registros[3674]= 3'b100;  
registros[3675]= 3'b000;  
registros[3676]= 3'b000;  
registros[3677]= 3'b000;  
registros[3678]= 3'b000;  
registros[3679]= 3'b000;  
registros[3680]= 3'b000;  
registros[3681]= 3'b000;  
registros[3682]= 3'b000;  
registros[3683]= 3'b000;  
registros[3684]= 3'b000;  
registros[3685]= 3'b000;  
registros[3686]= 3'b000;  
registros[3687]= 3'b000;  
registros[3688]= 3'b000;  
registros[3689]= 3'b000;  
registros[3690]= 3'b000;  
registros[3691]= 3'b111;  
registros[3692]= 3'b111;  
registros[3693]= 3'b111;  
registros[3694]= 3'b111;  
registros[3695]= 3'b111;  
registros[3696]= 3'b111;  
registros[3697]= 3'b111;  
registros[3698]= 3'b111;  
registros[3699]= 3'b111;  
registros[3700]= 3'b111;  
registros[3701]= 3'b111;  
registros[3702]= 3'b111;  
registros[3703]= 3'b111;  
registros[3704]= 3'b111;  
registros[3705]= 3'b111;  
registros[3706]= 3'b111;  
registros[3707]= 3'b111;  
registros[3708]= 3'b111;  
registros[3709]= 3'b111;  
registros[3710]= 3'b111;  
registros[3711]= 3'b111;  
registros[3712]= 3'b111;  
registros[3713]= 3'b111;  
registros[3714]= 3'b111;  
registros[3715]= 3'b111;  
registros[3716]= 3'b111;  
registros[3717]= 3'b111;  
registros[3718]= 3'b111;  
registros[3719]= 3'b111;  
registros[3720]= 3'b111;  
registros[3721]= 3'b111;  
registros[3722]= 3'b111;  
registros[3723]= 3'b000;  
registros[3724]= 3'b000;  
registros[3725]= 3'b000;  
registros[3726]= 3'b000;  
registros[3727]= 3'b100;  
registros[3728]= 3'b100;  
registros[3729]= 3'b100;  
registros[3730]= 3'b000;  
registros[3731]= 3'b000;  
registros[3732]= 3'b100;  
registros[3733]= 3'b100;  
registros[3734]= 3'b100;  
registros[3735]= 3'b100;  
registros[3736]= 3'b100;  
registros[3737]= 3'b100;  
registros[3738]= 3'b000;  
registros[3739]= 3'b000;  
registros[3740]= 3'b000;  
registros[3741]= 3'b000;  
registros[3742]= 3'b000;  
registros[3743]= 3'b000;  
registros[3744]= 3'b000;  
registros[3745]= 3'b000;  
registros[3746]= 3'b000;  
registros[3747]= 3'b000;  
registros[3748]= 3'b000;  
registros[3749]= 3'b000;  
registros[3750]= 3'b000;  
registros[3751]= 3'b000;  
registros[3752]= 3'b000;  
registros[3753]= 3'b111;  
registros[3754]= 3'b111;  
registros[3755]= 3'b111;  
registros[3756]= 3'b111;  
registros[3757]= 3'b111;  
registros[3758]= 3'b111;  
registros[3759]= 3'b111;  
registros[3760]= 3'b111;  
registros[3761]= 3'b111;  
registros[3762]= 3'b111;  
registros[3763]= 3'b111;  
registros[3764]= 3'b111;  
registros[3765]= 3'b111;  
registros[3766]= 3'b111;  
registros[3767]= 3'b111;  
registros[3768]= 3'b111;  
registros[3769]= 3'b111;  
registros[3770]= 3'b111;  
registros[3771]= 3'b111;  
registros[3772]= 3'b111;  
registros[3773]= 3'b111;  
registros[3774]= 3'b111;  
registros[3775]= 3'b111;  
registros[3776]= 3'b111;  
registros[3777]= 3'b111;  
registros[3778]= 3'b111;  
registros[3779]= 3'b111;  
registros[3780]= 3'b111;  
registros[3781]= 3'b111;  
registros[3782]= 3'b111;  
registros[3783]= 3'b111;  
registros[3784]= 3'b111;  
registros[3785]= 3'b111;  
registros[3786]= 3'b111;  
registros[3787]= 3'b111;  
registros[3788]= 3'b111;  
registros[3789]= 3'b111;  
registros[3790]= 3'b111;  
registros[3791]= 3'b111;  
registros[3792]= 3'b111;  
registros[3793]= 3'b000;  
registros[3794]= 3'b000;  
registros[3795]= 3'b100;  
registros[3796]= 3'b100;  
registros[3797]= 3'b100;  
registros[3798]= 3'b100;  
registros[3799]= 3'b100;  
registros[3800]= 3'b100;  
registros[3801]= 3'b000;  
registros[3802]= 3'b000;  
registros[3803]= 3'b000;  
registros[3804]= 3'b000;  
registros[3805]= 3'b000;  
registros[3806]= 3'b000;  
registros[3807]= 3'b000;  
registros[3808]= 3'b000;  
registros[3809]= 3'b000;  
registros[3810]= 3'b000;  
registros[3811]= 3'b000;  
registros[3812]= 3'b000;  
registros[3813]= 3'b000;  
registros[3814]= 3'b111;  
registros[3815]= 3'b111;  
registros[3816]= 3'b111;  
registros[3817]= 3'b111;  
registros[3818]= 3'b111;  
registros[3819]= 3'b111;  
registros[3820]= 3'b111;  
registros[3821]= 3'b111;  
registros[3822]= 3'b111;  
registros[3823]= 3'b111;  
registros[3824]= 3'b111;  
registros[3825]= 3'b111;  
registros[3826]= 3'b111;  
registros[3827]= 3'b111;  
registros[3828]= 3'b111;  
registros[3829]= 3'b111;  
registros[3830]= 3'b111;  
registros[3831]= 3'b111;  
registros[3832]= 3'b111;  
registros[3833]= 3'b111;  
registros[3834]= 3'b111;  
registros[3835]= 3'b111;  
registros[3836]= 3'b111;  
registros[3837]= 3'b111;  
registros[3838]= 3'b111;  
registros[3839]= 3'b111;  
registros[3840]= 3'b111;  
registros[3841]= 3'b111;  
registros[3842]= 3'b111;  
registros[3843]= 3'b111;  
registros[3844]= 3'b111;  
registros[3845]= 3'b111;  
registros[3846]= 3'b111;  
registros[3847]= 3'b111;  
registros[3848]= 3'b111;  
registros[3849]= 3'b111;  
registros[3850]= 3'b111;  
registros[3851]= 3'b111;  
registros[3852]= 3'b111;  
registros[3853]= 3'b111;  
registros[3854]= 3'b111;  
registros[3855]= 3'b111;  
registros[3856]= 3'b111;  
registros[3857]= 3'b111;  
registros[3858]= 3'b000;  
registros[3859]= 3'b000;  
registros[3860]= 3'b000;  
registros[3861]= 3'b100;  
registros[3862]= 3'b100;  
registros[3863]= 3'b100;  
registros[3864]= 3'b000;  
registros[3865]= 3'b000;  
registros[3866]= 3'b000;  
registros[3867]= 3'b000;  
registros[3868]= 3'b000;  
registros[3869]= 3'b000;  
registros[3870]= 3'b000;  
registros[3871]= 3'b000;  
registros[3872]= 3'b000;  
registros[3873]= 3'b000;  
registros[3874]= 3'b000;  
registros[3875]= 3'b000;  
registros[3876]= 3'b000;  
registros[3877]= 3'b111;  
registros[3878]= 3'b111;  
registros[3879]= 3'b111;  
registros[3880]= 3'b111;  
registros[3881]= 3'b111;  
registros[3882]= 3'b111;  
registros[3883]= 3'b111;  
registros[3884]= 3'b111;  
registros[3885]= 3'b111;  
registros[3886]= 3'b111;  
registros[3887]= 3'b111;  
registros[3888]= 3'b111;  
registros[3889]= 3'b111;  
registros[3890]= 3'b111;  
registros[3891]= 3'b111;  
registros[3892]= 3'b111;  
registros[3893]= 3'b111;  
registros[3894]= 3'b111;  
registros[3895]= 3'b111;  
registros[3896]= 3'b111;  
registros[3897]= 3'b111;  
registros[3898]= 3'b111;  
registros[3899]= 3'b111;  
registros[3900]= 3'b111;  
registros[3901]= 3'b111;  
registros[3902]= 3'b111;  
registros[3903]= 3'b111;  
registros[3904]= 3'b111;  
registros[3905]= 3'b111;  
registros[3906]= 3'b111;  
registros[3907]= 3'b111;  
registros[3908]= 3'b111;  
registros[3909]= 3'b111;  
registros[3910]= 3'b111;  
registros[3911]= 3'b111;  
registros[3912]= 3'b111;  
registros[3913]= 3'b111;  
registros[3914]= 3'b111;  
registros[3915]= 3'b111;  
registros[3916]= 3'b111;  
registros[3917]= 3'b111;  
registros[3918]= 3'b111;  
registros[3919]= 3'b111;  
registros[3920]= 3'b111;  
registros[3921]= 3'b111;  
registros[3922]= 3'b111;  
registros[3923]= 3'b111;  
registros[3924]= 3'b111;  
registros[3925]= 3'b000;  
registros[3926]= 3'b000;  
registros[3927]= 3'b000;  
registros[3928]= 3'b000;  
registros[3929]= 3'b000;  
registros[3930]= 3'b000;  
registros[3931]= 3'b000;  
registros[3932]= 3'b000;  
registros[3933]= 3'b000;  
registros[3934]= 3'b000;  
registros[3935]= 3'b000;  
registros[3936]= 3'b000;  
registros[3937]= 3'b000;  
registros[3938]= 3'b000;  
registros[3939]= 3'b000;  
registros[3940]= 3'b111;  
registros[3941]= 3'b111;  
registros[3942]= 3'b111;  
registros[3943]= 3'b111;  
registros[3944]= 3'b111;  
registros[3945]= 3'b111;  
registros[3946]= 3'b111;  
registros[3947]= 3'b111;  
registros[3948]= 3'b111;  
registros[3949]= 3'b111;  
registros[3950]= 3'b111;  
registros[3951]= 3'b111;  
registros[3952]= 3'b111;  
registros[3953]= 3'b111;  
registros[3954]= 3'b111;  
registros[3955]= 3'b111;  
registros[3956]= 3'b111;  
registros[3957]= 3'b111;  
registros[3958]= 3'b111;  
registros[3959]= 3'b111;  
registros[3960]= 3'b111;  
registros[3961]= 3'b111;  
registros[3962]= 3'b111;  
registros[3963]= 3'b111;  
registros[3964]= 3'b111;  
registros[3965]= 3'b111;  
registros[3966]= 3'b111;  
registros[3967]= 3'b111;  
registros[3968]= 3'b111;  
registros[3969]= 3'b111;  
registros[3970]= 3'b111;  
registros[3971]= 3'b111;  
registros[3972]= 3'b111;  
registros[3973]= 3'b111;  
registros[3974]= 3'b111;  
registros[3975]= 3'b111;  
registros[3976]= 3'b111;  
registros[3977]= 3'b111;  
registros[3978]= 3'b111;  
registros[3979]= 3'b111;  
registros[3980]= 3'b111;  
registros[3981]= 3'b111;  
registros[3982]= 3'b111;  
registros[3983]= 3'b111;  
registros[3984]= 3'b111;  
registros[3985]= 3'b111;  
registros[3986]= 3'b111;  
registros[3987]= 3'b111;  
registros[3988]= 3'b111;  
registros[3989]= 3'b111;  
registros[3990]= 3'b111;  
registros[3991]= 3'b000;  
registros[3992]= 3'b000;  
registros[3993]= 3'b000;  
registros[3994]= 3'b000;  
registros[3995]= 3'b000;  
registros[3996]= 3'b000;  
registros[3997]= 3'b000;  
registros[3998]= 3'b000;  
registros[3999]= 3'b000;  
registros[4000]= 3'b000;  
registros[4001]= 3'b000;  
registros[4002]= 3'b111;  
registros[4003]= 3'b111;  
registros[4004]= 3'b111;  
registros[4005]= 3'b111;  
registros[4006]= 3'b111;  
registros[4007]= 3'b111;  
registros[4008]= 3'b111;  
registros[4009]= 3'b111;  
registros[4010]= 3'b111;  
registros[4011]= 3'b111;  
registros[4012]= 3'b111;  
registros[4013]= 3'b111;  
registros[4014]= 3'b111;  
registros[4015]= 3'b111;  
registros[4016]= 3'b111;  
registros[4017]= 3'b111;  
registros[4018]= 3'b111;  
registros[4019]= 3'b111;  
registros[4020]= 3'b111;  
registros[4021]= 3'b111;  
registros[4022]= 3'b111;  
registros[4023]= 3'b111;  
registros[4024]= 3'b111;  
registros[4025]= 3'b111;  
registros[4026]= 3'b111;  
registros[4027]= 3'b111;  
registros[4028]= 3'b111;  
registros[4029]= 3'b111;  
registros[4030]= 3'b111;  
registros[4031]= 3'b111;  
registros[4032]= 3'b111;  
registros[4033]= 3'b111;  
registros[4034]= 3'b111;  
registros[4035]= 3'b111;  
registros[4036]= 3'b111;  
registros[4037]= 3'b111;  
registros[4038]= 3'b111;  
registros[4039]= 3'b111;  
registros[4040]= 3'b111;  
registros[4041]= 3'b111;  
registros[4042]= 3'b111;  
registros[4043]= 3'b111;  
registros[4044]= 3'b111;  
registros[4045]= 3'b111;  
registros[4046]= 3'b111;  
registros[4047]= 3'b111;  
registros[4048]= 3'b111;  
registros[4049]= 3'b111;  
registros[4050]= 3'b111;  
registros[4051]= 3'b111;  
registros[4052]= 3'b111;  
registros[4053]= 3'b111;  
registros[4054]= 3'b111;  
registros[4055]= 3'b111;  
registros[4056]= 3'b111;  
registros[4057]= 3'b111;  
registros[4058]= 3'b000;  
registros[4059]= 3'b000;  
registros[4060]= 3'b000;  
registros[4061]= 3'b000;  
registros[4062]= 3'b000;  
registros[4063]= 3'b000;  
registros[4064]= 3'b111;  
registros[4065]= 3'b111;  
registros[4066]= 3'b111;  
registros[4067]= 3'b111;  
registros[4068]= 3'b111;  
registros[4069]= 3'b111;  
registros[4070]= 3'b111;  
registros[4071]= 3'b111;  
registros[4072]= 3'b111;  
registros[4073]= 3'b111;  
registros[4074]= 3'b111;  
registros[4075]= 3'b111;  
registros[4076]= 3'b111;  
registros[4077]= 3'b111;  
registros[4078]= 3'b111;  
registros[4079]= 3'b111;  
registros[4080]= 3'b111;  
registros[4081]= 3'b111;  
registros[4082]= 3'b111;  
registros[4083]= 3'b111;  
registros[4084]= 3'b111;  
registros[4085]= 3'b111;  
registros[4086]= 3'b111;  
registros[4087]= 3'b111;  
registros[4088]= 3'b111;  
registros[4089]= 3'b111;  
registros[4090]= 3'b111;  
registros[4091]= 3'b111;  
registros[4092]= 3'b111;  
registros[4093]= 3'b111;  
registros[4094]= 3'b111;  
registros[4095]= 3'b111;  
end

always @(posedge clk) begin
	if(hcount>10'd550 || hcount<10'd190)
		w_rgb = 4'b1000;
	else if (hcount>=origen_x && hcount<(origen_x+tamano) && vcount<(y_tamano + origen_y) && vcount>= origen_y) begin
		w_rgb = {1'b0,registros[lectura]};
	end
	else begin
		w_rgb = 4'b1000;
	end
end

assign rgb_out = w_rgb;
assign lectura = (vcount - origen_y)*tamano + (hcount - origen_x);

endmodule
